
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"fc",x"f5",x"c2",x"87"),
    12 => (x"48",x"c0",x"c8",x"4e"),
    13 => (x"d5",x"c1",x"28",x"c2"),
    14 => (x"ea",x"d6",x"e5",x"ea"),
    15 => (x"c1",x"46",x"71",x"49"),
    16 => (x"87",x"f9",x"01",x"88"),
    17 => (x"49",x"fc",x"f5",x"c2"),
    18 => (x"48",x"c4",x"e3",x"c2"),
    19 => (x"03",x"89",x"d0",x"89"),
    20 => (x"40",x"40",x"40",x"c0"),
    21 => (x"d0",x"87",x"f6",x"40"),
    22 => (x"50",x"c0",x"05",x"81"),
    23 => (x"f9",x"05",x"89",x"c1"),
    24 => (x"c4",x"e3",x"c2",x"87"),
    25 => (x"c0",x"e3",x"c2",x"4d"),
    26 => (x"02",x"ad",x"74",x"4c"),
    27 => (x"0f",x"24",x"87",x"c4"),
    28 => (x"e8",x"c1",x"87",x"f7"),
    29 => (x"e3",x"c2",x"87",x"c6"),
    30 => (x"e3",x"c2",x"4d",x"c4"),
    31 => (x"ad",x"74",x"4c",x"c4"),
    32 => (x"c4",x"87",x"c6",x"02"),
    33 => (x"f5",x"0f",x"6c",x"8c"),
    34 => (x"87",x"fd",x"00",x"87"),
    35 => (x"71",x"86",x"fc",x"1e"),
    36 => (x"49",x"c0",x"ff",x"4a"),
    37 => (x"c0",x"c4",x"48",x"69"),
    38 => (x"48",x"7e",x"70",x"98"),
    39 => (x"87",x"f4",x"02",x"98"),
    40 => (x"fc",x"48",x"79",x"72"),
    41 => (x"0e",x"4f",x"26",x"8e"),
    42 => (x"0e",x"5c",x"5b",x"5e"),
    43 => (x"4c",x"c0",x"4b",x"71"),
    44 => (x"02",x"9a",x"4a",x"13"),
    45 => (x"49",x"72",x"87",x"cd"),
    46 => (x"c1",x"87",x"d1",x"ff"),
    47 => (x"9a",x"4a",x"13",x"84"),
    48 => (x"74",x"87",x"f3",x"05"),
    49 => (x"26",x"4c",x"26",x"48"),
    50 => (x"1e",x"4f",x"26",x"4b"),
    51 => (x"1e",x"73",x"1e",x"72"),
    52 => (x"02",x"11",x"48",x"12"),
    53 => (x"c3",x"4b",x"87",x"ca"),
    54 => (x"73",x"9b",x"98",x"df"),
    55 => (x"87",x"f0",x"02",x"88"),
    56 => (x"4a",x"26",x"4b",x"26"),
    57 => (x"73",x"1e",x"4f",x"26"),
    58 => (x"c1",x"1e",x"72",x"1e"),
    59 => (x"87",x"ca",x"04",x"8b"),
    60 => (x"02",x"11",x"48",x"12"),
    61 => (x"02",x"88",x"87",x"c4"),
    62 => (x"4a",x"26",x"87",x"f1"),
    63 => (x"4f",x"26",x"4b",x"26"),
    64 => (x"73",x"1e",x"74",x"1e"),
    65 => (x"c1",x"1e",x"72",x"1e"),
    66 => (x"87",x"d0",x"04",x"8b"),
    67 => (x"02",x"11",x"48",x"12"),
    68 => (x"c3",x"4c",x"87",x"ca"),
    69 => (x"74",x"9c",x"98",x"df"),
    70 => (x"87",x"eb",x"02",x"88"),
    71 => (x"4b",x"26",x"4a",x"26"),
    72 => (x"4f",x"26",x"4c",x"26"),
    73 => (x"81",x"48",x"73",x"1e"),
    74 => (x"c5",x"02",x"a9",x"73"),
    75 => (x"05",x"53",x"12",x"87"),
    76 => (x"4f",x"26",x"87",x"f6"),
    77 => (x"71",x"1e",x"73",x"1e"),
    78 => (x"4b",x"66",x"c8",x"4a"),
    79 => (x"71",x"8b",x"c1",x"49"),
    80 => (x"87",x"cf",x"02",x"99"),
    81 => (x"d4",x"ff",x"48",x"12"),
    82 => (x"49",x"73",x"78",x"08"),
    83 => (x"99",x"71",x"8b",x"c1"),
    84 => (x"26",x"87",x"f1",x"05"),
    85 => (x"0e",x"4f",x"26",x"4b"),
    86 => (x"0e",x"5c",x"5b",x"5e"),
    87 => (x"d4",x"ff",x"4a",x"71"),
    88 => (x"4b",x"66",x"cc",x"4c"),
    89 => (x"71",x"8b",x"c1",x"49"),
    90 => (x"87",x"ce",x"02",x"99"),
    91 => (x"6c",x"7c",x"ff",x"c3"),
    92 => (x"c1",x"49",x"73",x"52"),
    93 => (x"05",x"99",x"71",x"8b"),
    94 => (x"4c",x"26",x"87",x"f2"),
    95 => (x"4f",x"26",x"4b",x"26"),
    96 => (x"ff",x"1e",x"73",x"1e"),
    97 => (x"ff",x"c3",x"4b",x"d4"),
    98 => (x"c3",x"4a",x"6b",x"7b"),
    99 => (x"49",x"6b",x"7b",x"ff"),
   100 => (x"b1",x"72",x"32",x"c8"),
   101 => (x"6b",x"7b",x"ff",x"c3"),
   102 => (x"71",x"31",x"c8",x"4a"),
   103 => (x"7b",x"ff",x"c3",x"b2"),
   104 => (x"32",x"c8",x"49",x"6b"),
   105 => (x"48",x"71",x"b1",x"72"),
   106 => (x"4f",x"26",x"4b",x"26"),
   107 => (x"5c",x"5b",x"5e",x"0e"),
   108 => (x"4d",x"71",x"0e",x"5d"),
   109 => (x"75",x"4c",x"d4",x"ff"),
   110 => (x"98",x"ff",x"c3",x"48"),
   111 => (x"e3",x"c2",x"7c",x"70"),
   112 => (x"c8",x"05",x"bf",x"c4"),
   113 => (x"48",x"66",x"d0",x"87"),
   114 => (x"a6",x"d4",x"30",x"c9"),
   115 => (x"49",x"66",x"d0",x"58"),
   116 => (x"48",x"71",x"29",x"d8"),
   117 => (x"70",x"98",x"ff",x"c3"),
   118 => (x"49",x"66",x"d0",x"7c"),
   119 => (x"48",x"71",x"29",x"d0"),
   120 => (x"70",x"98",x"ff",x"c3"),
   121 => (x"49",x"66",x"d0",x"7c"),
   122 => (x"48",x"71",x"29",x"c8"),
   123 => (x"70",x"98",x"ff",x"c3"),
   124 => (x"48",x"66",x"d0",x"7c"),
   125 => (x"70",x"98",x"ff",x"c3"),
   126 => (x"d0",x"49",x"75",x"7c"),
   127 => (x"c3",x"48",x"71",x"29"),
   128 => (x"7c",x"70",x"98",x"ff"),
   129 => (x"f0",x"c9",x"4b",x"6c"),
   130 => (x"ff",x"c3",x"4a",x"ff"),
   131 => (x"87",x"cf",x"05",x"ab"),
   132 => (x"6c",x"7c",x"71",x"49"),
   133 => (x"02",x"8a",x"c1",x"4b"),
   134 => (x"ab",x"71",x"87",x"c5"),
   135 => (x"73",x"87",x"f2",x"02"),
   136 => (x"26",x"4d",x"26",x"48"),
   137 => (x"26",x"4b",x"26",x"4c"),
   138 => (x"49",x"c0",x"1e",x"4f"),
   139 => (x"c3",x"48",x"d4",x"ff"),
   140 => (x"81",x"c1",x"78",x"ff"),
   141 => (x"a9",x"b7",x"c8",x"c3"),
   142 => (x"26",x"87",x"f1",x"04"),
   143 => (x"5b",x"5e",x"0e",x"4f"),
   144 => (x"c0",x"0e",x"5d",x"5c"),
   145 => (x"f7",x"c1",x"f0",x"ff"),
   146 => (x"c0",x"c0",x"c1",x"4d"),
   147 => (x"4b",x"c0",x"c0",x"c0"),
   148 => (x"c4",x"87",x"d6",x"ff"),
   149 => (x"c0",x"4c",x"df",x"f8"),
   150 => (x"fd",x"49",x"75",x"1e"),
   151 => (x"86",x"c4",x"87",x"ce"),
   152 => (x"c0",x"05",x"a8",x"c1"),
   153 => (x"d4",x"ff",x"87",x"e5"),
   154 => (x"78",x"ff",x"c3",x"48"),
   155 => (x"e1",x"c0",x"1e",x"73"),
   156 => (x"49",x"e9",x"c1",x"f0"),
   157 => (x"c4",x"87",x"f5",x"fc"),
   158 => (x"05",x"98",x"70",x"86"),
   159 => (x"d4",x"ff",x"87",x"ca"),
   160 => (x"78",x"ff",x"c3",x"48"),
   161 => (x"87",x"cb",x"48",x"c1"),
   162 => (x"c1",x"87",x"de",x"fe"),
   163 => (x"c6",x"ff",x"05",x"8c"),
   164 => (x"26",x"48",x"c0",x"87"),
   165 => (x"26",x"4c",x"26",x"4d"),
   166 => (x"0e",x"4f",x"26",x"4b"),
   167 => (x"0e",x"5c",x"5b",x"5e"),
   168 => (x"c1",x"f0",x"ff",x"c0"),
   169 => (x"d4",x"ff",x"4c",x"c1"),
   170 => (x"78",x"ff",x"c3",x"48"),
   171 => (x"f7",x"49",x"e0",x"cb"),
   172 => (x"4b",x"d3",x"87",x"f5"),
   173 => (x"49",x"74",x"1e",x"c0"),
   174 => (x"c4",x"87",x"f1",x"fb"),
   175 => (x"05",x"98",x"70",x"86"),
   176 => (x"d4",x"ff",x"87",x"ca"),
   177 => (x"78",x"ff",x"c3",x"48"),
   178 => (x"87",x"cb",x"48",x"c1"),
   179 => (x"c1",x"87",x"da",x"fd"),
   180 => (x"df",x"ff",x"05",x"8b"),
   181 => (x"26",x"48",x"c0",x"87"),
   182 => (x"26",x"4b",x"26",x"4c"),
   183 => (x"00",x"00",x"00",x"4f"),
   184 => (x"00",x"44",x"4d",x"43"),
   185 => (x"5c",x"5b",x"5e",x"0e"),
   186 => (x"ff",x"c3",x"0e",x"5d"),
   187 => (x"4b",x"d4",x"ff",x"4d"),
   188 => (x"c6",x"87",x"f6",x"fc"),
   189 => (x"e1",x"c0",x"1e",x"ea"),
   190 => (x"49",x"c8",x"c1",x"f0"),
   191 => (x"c4",x"87",x"ed",x"fa"),
   192 => (x"02",x"a8",x"c1",x"86"),
   193 => (x"d2",x"fe",x"87",x"c8"),
   194 => (x"c1",x"48",x"c0",x"87"),
   195 => (x"ef",x"f9",x"87",x"e8"),
   196 => (x"cf",x"49",x"70",x"87"),
   197 => (x"c6",x"99",x"ff",x"ff"),
   198 => (x"c8",x"02",x"a9",x"ea"),
   199 => (x"87",x"fb",x"fd",x"87"),
   200 => (x"d1",x"c1",x"48",x"c0"),
   201 => (x"c0",x"7b",x"75",x"87"),
   202 => (x"d0",x"fc",x"4c",x"f1"),
   203 => (x"02",x"98",x"70",x"87"),
   204 => (x"c0",x"87",x"ec",x"c0"),
   205 => (x"f0",x"ff",x"c0",x"1e"),
   206 => (x"f9",x"49",x"fa",x"c1"),
   207 => (x"86",x"c4",x"87",x"ee"),
   208 => (x"da",x"05",x"98",x"70"),
   209 => (x"6b",x"7b",x"75",x"87"),
   210 => (x"75",x"7b",x"75",x"49"),
   211 => (x"75",x"7b",x"75",x"7b"),
   212 => (x"99",x"c0",x"c1",x"7b"),
   213 => (x"c1",x"87",x"c4",x"02"),
   214 => (x"c0",x"87",x"db",x"48"),
   215 => (x"c2",x"87",x"d7",x"48"),
   216 => (x"87",x"ca",x"05",x"ac"),
   217 => (x"f4",x"49",x"c0",x"ce"),
   218 => (x"48",x"c0",x"87",x"fd"),
   219 => (x"8c",x"c1",x"87",x"c8"),
   220 => (x"87",x"f6",x"fe",x"05"),
   221 => (x"4d",x"26",x"48",x"c0"),
   222 => (x"4b",x"26",x"4c",x"26"),
   223 => (x"00",x"00",x"4f",x"26"),
   224 => (x"43",x"48",x"44",x"53"),
   225 => (x"69",x"61",x"66",x"20"),
   226 => (x"00",x"0a",x"21",x"6c"),
   227 => (x"5c",x"5b",x"5e",x"0e"),
   228 => (x"d0",x"ff",x"0e",x"5d"),
   229 => (x"d0",x"e5",x"c0",x"4d"),
   230 => (x"c2",x"4c",x"c0",x"c1"),
   231 => (x"c1",x"48",x"c4",x"e3"),
   232 => (x"49",x"d8",x"d0",x"78"),
   233 => (x"c7",x"87",x"c0",x"f4"),
   234 => (x"f9",x"7d",x"c2",x"4b"),
   235 => (x"7d",x"c3",x"87",x"fb"),
   236 => (x"49",x"74",x"1e",x"c0"),
   237 => (x"c4",x"87",x"f5",x"f7"),
   238 => (x"05",x"a8",x"c1",x"86"),
   239 => (x"c2",x"4b",x"87",x"c1"),
   240 => (x"87",x"cb",x"05",x"ab"),
   241 => (x"f3",x"49",x"d0",x"d0"),
   242 => (x"48",x"c0",x"87",x"dd"),
   243 => (x"c1",x"87",x"f6",x"c0"),
   244 => (x"d4",x"ff",x"05",x"8b"),
   245 => (x"87",x"cc",x"fc",x"87"),
   246 => (x"58",x"c8",x"e3",x"c2"),
   247 => (x"cd",x"05",x"98",x"70"),
   248 => (x"c0",x"1e",x"c1",x"87"),
   249 => (x"d0",x"c1",x"f0",x"ff"),
   250 => (x"87",x"c0",x"f7",x"49"),
   251 => (x"d4",x"ff",x"86",x"c4"),
   252 => (x"78",x"ff",x"c3",x"48"),
   253 => (x"c2",x"87",x"cc",x"c5"),
   254 => (x"c2",x"58",x"cc",x"e3"),
   255 => (x"48",x"d4",x"ff",x"7d"),
   256 => (x"c1",x"78",x"ff",x"c3"),
   257 => (x"26",x"4d",x"26",x"48"),
   258 => (x"26",x"4b",x"26",x"4c"),
   259 => (x"00",x"00",x"00",x"4f"),
   260 => (x"52",x"52",x"45",x"49"),
   261 => (x"00",x"00",x"00",x"00"),
   262 => (x"00",x"49",x"50",x"53"),
   263 => (x"5c",x"5b",x"5e",x"0e"),
   264 => (x"4d",x"71",x"0e",x"5d"),
   265 => (x"ff",x"4c",x"ff",x"c3"),
   266 => (x"7b",x"74",x"4b",x"d4"),
   267 => (x"c4",x"48",x"d0",x"ff"),
   268 => (x"7b",x"74",x"78",x"c3"),
   269 => (x"ff",x"c0",x"1e",x"75"),
   270 => (x"49",x"d8",x"c1",x"f0"),
   271 => (x"c4",x"87",x"ed",x"f5"),
   272 => (x"02",x"98",x"70",x"86"),
   273 => (x"c8",x"d2",x"87",x"cb"),
   274 => (x"87",x"db",x"f1",x"49"),
   275 => (x"ee",x"c0",x"48",x"c1"),
   276 => (x"c3",x"7b",x"74",x"87"),
   277 => (x"c0",x"c8",x"7b",x"fe"),
   278 => (x"49",x"66",x"d4",x"1e"),
   279 => (x"c4",x"87",x"d5",x"f3"),
   280 => (x"74",x"7b",x"74",x"86"),
   281 => (x"d8",x"7b",x"74",x"7b"),
   282 => (x"74",x"4a",x"e0",x"da"),
   283 => (x"c5",x"05",x"6b",x"7b"),
   284 => (x"05",x"8a",x"c1",x"87"),
   285 => (x"7b",x"74",x"87",x"f5"),
   286 => (x"c2",x"48",x"d0",x"ff"),
   287 => (x"26",x"48",x"c0",x"78"),
   288 => (x"26",x"4c",x"26",x"4d"),
   289 => (x"00",x"4f",x"26",x"4b"),
   290 => (x"74",x"69",x"72",x"57"),
   291 => (x"61",x"66",x"20",x"65"),
   292 => (x"64",x"65",x"6c",x"69"),
   293 => (x"5e",x"0e",x"00",x"0a"),
   294 => (x"0e",x"5d",x"5c",x"5b"),
   295 => (x"4b",x"71",x"86",x"fc"),
   296 => (x"c0",x"4c",x"d4",x"ff"),
   297 => (x"cd",x"ee",x"c5",x"7e"),
   298 => (x"ff",x"c3",x"4a",x"df"),
   299 => (x"c3",x"48",x"6c",x"7c"),
   300 => (x"c0",x"05",x"a8",x"fe"),
   301 => (x"4d",x"74",x"87",x"f8"),
   302 => (x"cc",x"02",x"9b",x"73"),
   303 => (x"1e",x"66",x"d4",x"87"),
   304 => (x"d2",x"f2",x"49",x"73"),
   305 => (x"d4",x"86",x"c4",x"87"),
   306 => (x"48",x"d0",x"ff",x"87"),
   307 => (x"d4",x"78",x"d1",x"c4"),
   308 => (x"ff",x"c3",x"4a",x"66"),
   309 => (x"05",x"8a",x"c1",x"7d"),
   310 => (x"a6",x"d8",x"87",x"f8"),
   311 => (x"7c",x"ff",x"c3",x"5a"),
   312 => (x"05",x"9b",x"73",x"7c"),
   313 => (x"d0",x"ff",x"87",x"c5"),
   314 => (x"c1",x"78",x"d0",x"48"),
   315 => (x"8a",x"c1",x"7e",x"4a"),
   316 => (x"87",x"f6",x"fe",x"05"),
   317 => (x"8e",x"fc",x"48",x"6e"),
   318 => (x"4c",x"26",x"4d",x"26"),
   319 => (x"4f",x"26",x"4b",x"26"),
   320 => (x"71",x"1e",x"73",x"1e"),
   321 => (x"ff",x"4b",x"c0",x"4a"),
   322 => (x"ff",x"c3",x"48",x"d4"),
   323 => (x"48",x"d0",x"ff",x"78"),
   324 => (x"ff",x"78",x"c3",x"c4"),
   325 => (x"ff",x"c3",x"48",x"d4"),
   326 => (x"c0",x"1e",x"72",x"78"),
   327 => (x"d1",x"c1",x"f0",x"ff"),
   328 => (x"87",x"c8",x"f2",x"49"),
   329 => (x"98",x"70",x"86",x"c4"),
   330 => (x"c8",x"87",x"d2",x"05"),
   331 => (x"66",x"cc",x"1e",x"c0"),
   332 => (x"87",x"e2",x"fd",x"49"),
   333 => (x"4b",x"70",x"86",x"c4"),
   334 => (x"c2",x"48",x"d0",x"ff"),
   335 => (x"26",x"48",x"73",x"78"),
   336 => (x"0e",x"4f",x"26",x"4b"),
   337 => (x"5d",x"5c",x"5b",x"5e"),
   338 => (x"c0",x"1e",x"c0",x"0e"),
   339 => (x"c9",x"c1",x"f0",x"ff"),
   340 => (x"87",x"d8",x"f1",x"49"),
   341 => (x"e3",x"c2",x"1e",x"d2"),
   342 => (x"f9",x"fc",x"49",x"cc"),
   343 => (x"c0",x"86",x"c8",x"87"),
   344 => (x"d2",x"84",x"c1",x"4c"),
   345 => (x"f8",x"04",x"ac",x"b7"),
   346 => (x"cc",x"e3",x"c2",x"87"),
   347 => (x"c3",x"49",x"bf",x"97"),
   348 => (x"c0",x"c1",x"99",x"c0"),
   349 => (x"e7",x"c0",x"05",x"a9"),
   350 => (x"d3",x"e3",x"c2",x"87"),
   351 => (x"d0",x"49",x"bf",x"97"),
   352 => (x"d4",x"e3",x"c2",x"31"),
   353 => (x"c8",x"4a",x"bf",x"97"),
   354 => (x"c2",x"b1",x"72",x"32"),
   355 => (x"bf",x"97",x"d5",x"e3"),
   356 => (x"4c",x"71",x"b1",x"4a"),
   357 => (x"ff",x"ff",x"ff",x"cf"),
   358 => (x"ca",x"84",x"c1",x"9c"),
   359 => (x"87",x"e7",x"c1",x"34"),
   360 => (x"97",x"d5",x"e3",x"c2"),
   361 => (x"31",x"c1",x"49",x"bf"),
   362 => (x"e3",x"c2",x"99",x"c6"),
   363 => (x"4a",x"bf",x"97",x"d6"),
   364 => (x"72",x"2a",x"b7",x"c7"),
   365 => (x"d1",x"e3",x"c2",x"b1"),
   366 => (x"4d",x"4a",x"bf",x"97"),
   367 => (x"e3",x"c2",x"9d",x"cf"),
   368 => (x"4a",x"bf",x"97",x"d2"),
   369 => (x"32",x"ca",x"9a",x"c3"),
   370 => (x"97",x"d3",x"e3",x"c2"),
   371 => (x"33",x"c2",x"4b",x"bf"),
   372 => (x"e3",x"c2",x"b2",x"73"),
   373 => (x"4b",x"bf",x"97",x"d4"),
   374 => (x"c6",x"9b",x"c0",x"c3"),
   375 => (x"b2",x"73",x"2b",x"b7"),
   376 => (x"48",x"c1",x"81",x"c2"),
   377 => (x"49",x"70",x"30",x"71"),
   378 => (x"30",x"75",x"48",x"c1"),
   379 => (x"4c",x"72",x"4d",x"70"),
   380 => (x"94",x"71",x"84",x"c1"),
   381 => (x"ad",x"b7",x"c0",x"c8"),
   382 => (x"c1",x"87",x"cc",x"06"),
   383 => (x"c8",x"2d",x"b7",x"34"),
   384 => (x"01",x"ad",x"b7",x"c0"),
   385 => (x"74",x"87",x"f4",x"ff"),
   386 => (x"26",x"4d",x"26",x"48"),
   387 => (x"26",x"4b",x"26",x"4c"),
   388 => (x"5b",x"5e",x"0e",x"4f"),
   389 => (x"f8",x"0e",x"5d",x"5c"),
   390 => (x"f4",x"eb",x"c2",x"86"),
   391 => (x"c2",x"78",x"c0",x"48"),
   392 => (x"c0",x"1e",x"ec",x"e3"),
   393 => (x"87",x"d8",x"fb",x"49"),
   394 => (x"98",x"70",x"86",x"c4"),
   395 => (x"c0",x"87",x"c5",x"05"),
   396 => (x"87",x"c0",x"c9",x"48"),
   397 => (x"7e",x"c1",x"4d",x"c0"),
   398 => (x"bf",x"d8",x"f7",x"c0"),
   399 => (x"e2",x"e4",x"c2",x"49"),
   400 => (x"4b",x"c8",x"71",x"4a"),
   401 => (x"70",x"87",x"df",x"ea"),
   402 => (x"87",x"c2",x"05",x"98"),
   403 => (x"f7",x"c0",x"7e",x"c0"),
   404 => (x"c2",x"49",x"bf",x"d4"),
   405 => (x"71",x"4a",x"fe",x"e4"),
   406 => (x"c9",x"ea",x"4b",x"c8"),
   407 => (x"05",x"98",x"70",x"87"),
   408 => (x"7e",x"c0",x"87",x"c2"),
   409 => (x"fd",x"c0",x"02",x"6e"),
   410 => (x"f2",x"ea",x"c2",x"87"),
   411 => (x"eb",x"c2",x"4d",x"bf"),
   412 => (x"7e",x"bf",x"9f",x"ea"),
   413 => (x"ea",x"d6",x"c5",x"48"),
   414 => (x"87",x"c7",x"05",x"a8"),
   415 => (x"bf",x"f2",x"ea",x"c2"),
   416 => (x"6e",x"87",x"ce",x"4d"),
   417 => (x"d5",x"e9",x"ca",x"48"),
   418 => (x"87",x"c5",x"02",x"a8"),
   419 => (x"e3",x"c7",x"48",x"c0"),
   420 => (x"ec",x"e3",x"c2",x"87"),
   421 => (x"f9",x"49",x"75",x"1e"),
   422 => (x"86",x"c4",x"87",x"e6"),
   423 => (x"c5",x"05",x"98",x"70"),
   424 => (x"c7",x"48",x"c0",x"87"),
   425 => (x"f7",x"c0",x"87",x"ce"),
   426 => (x"c2",x"49",x"bf",x"d4"),
   427 => (x"71",x"4a",x"fe",x"e4"),
   428 => (x"f1",x"e8",x"4b",x"c8"),
   429 => (x"05",x"98",x"70",x"87"),
   430 => (x"eb",x"c2",x"87",x"c8"),
   431 => (x"78",x"c1",x"48",x"f4"),
   432 => (x"f7",x"c0",x"87",x"da"),
   433 => (x"c2",x"49",x"bf",x"d8"),
   434 => (x"71",x"4a",x"e2",x"e4"),
   435 => (x"d5",x"e8",x"4b",x"c8"),
   436 => (x"02",x"98",x"70",x"87"),
   437 => (x"c0",x"87",x"c5",x"c0"),
   438 => (x"87",x"d8",x"c6",x"48"),
   439 => (x"97",x"ea",x"eb",x"c2"),
   440 => (x"d5",x"c1",x"49",x"bf"),
   441 => (x"cd",x"c0",x"05",x"a9"),
   442 => (x"eb",x"eb",x"c2",x"87"),
   443 => (x"c2",x"49",x"bf",x"97"),
   444 => (x"c0",x"02",x"a9",x"ea"),
   445 => (x"48",x"c0",x"87",x"c5"),
   446 => (x"c2",x"87",x"f9",x"c5"),
   447 => (x"bf",x"97",x"ec",x"e3"),
   448 => (x"e9",x"c3",x"48",x"7e"),
   449 => (x"ce",x"c0",x"02",x"a8"),
   450 => (x"c3",x"48",x"6e",x"87"),
   451 => (x"c0",x"02",x"a8",x"eb"),
   452 => (x"48",x"c0",x"87",x"c5"),
   453 => (x"c2",x"87",x"dd",x"c5"),
   454 => (x"bf",x"97",x"f7",x"e3"),
   455 => (x"c0",x"05",x"99",x"49"),
   456 => (x"e3",x"c2",x"87",x"cc"),
   457 => (x"49",x"bf",x"97",x"f8"),
   458 => (x"c0",x"02",x"a9",x"c2"),
   459 => (x"48",x"c0",x"87",x"c5"),
   460 => (x"c2",x"87",x"c1",x"c5"),
   461 => (x"bf",x"97",x"f9",x"e3"),
   462 => (x"f0",x"eb",x"c2",x"48"),
   463 => (x"48",x"4c",x"70",x"58"),
   464 => (x"eb",x"c2",x"88",x"c1"),
   465 => (x"e3",x"c2",x"58",x"f4"),
   466 => (x"49",x"bf",x"97",x"fa"),
   467 => (x"e3",x"c2",x"81",x"75"),
   468 => (x"4a",x"bf",x"97",x"fb"),
   469 => (x"a1",x"72",x"32",x"c8"),
   470 => (x"c4",x"f0",x"c2",x"7e"),
   471 => (x"c2",x"78",x"6e",x"48"),
   472 => (x"bf",x"97",x"fc",x"e3"),
   473 => (x"58",x"a6",x"c8",x"48"),
   474 => (x"bf",x"f4",x"eb",x"c2"),
   475 => (x"87",x"cf",x"c2",x"02"),
   476 => (x"bf",x"d4",x"f7",x"c0"),
   477 => (x"fe",x"e4",x"c2",x"49"),
   478 => (x"4b",x"c8",x"71",x"4a"),
   479 => (x"70",x"87",x"e7",x"e5"),
   480 => (x"c5",x"c0",x"02",x"98"),
   481 => (x"c3",x"48",x"c0",x"87"),
   482 => (x"eb",x"c2",x"87",x"ea"),
   483 => (x"c2",x"4c",x"bf",x"ec"),
   484 => (x"c2",x"5c",x"d8",x"f0"),
   485 => (x"bf",x"97",x"d1",x"e4"),
   486 => (x"c2",x"31",x"c8",x"49"),
   487 => (x"bf",x"97",x"d0",x"e4"),
   488 => (x"c2",x"49",x"a1",x"4a"),
   489 => (x"bf",x"97",x"d2",x"e4"),
   490 => (x"72",x"32",x"d0",x"4a"),
   491 => (x"e4",x"c2",x"49",x"a1"),
   492 => (x"4a",x"bf",x"97",x"d3"),
   493 => (x"a1",x"72",x"32",x"d8"),
   494 => (x"91",x"66",x"c4",x"49"),
   495 => (x"bf",x"c4",x"f0",x"c2"),
   496 => (x"cc",x"f0",x"c2",x"81"),
   497 => (x"d9",x"e4",x"c2",x"59"),
   498 => (x"c8",x"4a",x"bf",x"97"),
   499 => (x"d8",x"e4",x"c2",x"32"),
   500 => (x"a2",x"4b",x"bf",x"97"),
   501 => (x"da",x"e4",x"c2",x"4a"),
   502 => (x"d0",x"4b",x"bf",x"97"),
   503 => (x"4a",x"a2",x"73",x"33"),
   504 => (x"97",x"db",x"e4",x"c2"),
   505 => (x"9b",x"cf",x"4b",x"bf"),
   506 => (x"a2",x"73",x"33",x"d8"),
   507 => (x"d0",x"f0",x"c2",x"4a"),
   508 => (x"74",x"8a",x"c2",x"5a"),
   509 => (x"d0",x"f0",x"c2",x"92"),
   510 => (x"78",x"a1",x"72",x"48"),
   511 => (x"c2",x"87",x"c1",x"c1"),
   512 => (x"bf",x"97",x"fe",x"e3"),
   513 => (x"c2",x"31",x"c8",x"49"),
   514 => (x"bf",x"97",x"fd",x"e3"),
   515 => (x"c5",x"49",x"a1",x"4a"),
   516 => (x"81",x"ff",x"c7",x"31"),
   517 => (x"f0",x"c2",x"29",x"c9"),
   518 => (x"e4",x"c2",x"59",x"d8"),
   519 => (x"4a",x"bf",x"97",x"c3"),
   520 => (x"e4",x"c2",x"32",x"c8"),
   521 => (x"4b",x"bf",x"97",x"c2"),
   522 => (x"66",x"c4",x"4a",x"a2"),
   523 => (x"c2",x"82",x"6e",x"92"),
   524 => (x"c2",x"5a",x"d4",x"f0"),
   525 => (x"c0",x"48",x"cc",x"f0"),
   526 => (x"c8",x"f0",x"c2",x"78"),
   527 => (x"78",x"a1",x"72",x"48"),
   528 => (x"48",x"d8",x"f0",x"c2"),
   529 => (x"bf",x"cc",x"f0",x"c2"),
   530 => (x"dc",x"f0",x"c2",x"78"),
   531 => (x"d0",x"f0",x"c2",x"48"),
   532 => (x"eb",x"c2",x"78",x"bf"),
   533 => (x"c0",x"02",x"bf",x"f4"),
   534 => (x"48",x"74",x"87",x"c9"),
   535 => (x"7e",x"70",x"30",x"c4"),
   536 => (x"c2",x"87",x"c9",x"c0"),
   537 => (x"48",x"bf",x"d4",x"f0"),
   538 => (x"7e",x"70",x"30",x"c4"),
   539 => (x"48",x"f8",x"eb",x"c2"),
   540 => (x"48",x"c1",x"78",x"6e"),
   541 => (x"4d",x"26",x"8e",x"f8"),
   542 => (x"4b",x"26",x"4c",x"26"),
   543 => (x"5e",x"0e",x"4f",x"26"),
   544 => (x"0e",x"5d",x"5c",x"5b"),
   545 => (x"eb",x"c2",x"4a",x"71"),
   546 => (x"cb",x"02",x"bf",x"f4"),
   547 => (x"c7",x"4b",x"72",x"87"),
   548 => (x"c1",x"4d",x"72",x"2b"),
   549 => (x"87",x"c9",x"9d",x"ff"),
   550 => (x"2b",x"c8",x"4b",x"72"),
   551 => (x"ff",x"c3",x"4d",x"72"),
   552 => (x"c4",x"f0",x"c2",x"9d"),
   553 => (x"f7",x"c0",x"83",x"bf"),
   554 => (x"02",x"ab",x"bf",x"d0"),
   555 => (x"f7",x"c0",x"87",x"d9"),
   556 => (x"e3",x"c2",x"5b",x"d4"),
   557 => (x"49",x"73",x"1e",x"ec"),
   558 => (x"c4",x"87",x"c5",x"f1"),
   559 => (x"05",x"98",x"70",x"86"),
   560 => (x"48",x"c0",x"87",x"c5"),
   561 => (x"c2",x"87",x"e6",x"c0"),
   562 => (x"02",x"bf",x"f4",x"eb"),
   563 => (x"49",x"75",x"87",x"d2"),
   564 => (x"e3",x"c2",x"91",x"c4"),
   565 => (x"4c",x"69",x"81",x"ec"),
   566 => (x"ff",x"ff",x"ff",x"cf"),
   567 => (x"87",x"cb",x"9c",x"ff"),
   568 => (x"91",x"c2",x"49",x"75"),
   569 => (x"81",x"ec",x"e3",x"c2"),
   570 => (x"74",x"4c",x"69",x"9f"),
   571 => (x"26",x"4d",x"26",x"48"),
   572 => (x"26",x"4b",x"26",x"4c"),
   573 => (x"5b",x"5e",x"0e",x"4f"),
   574 => (x"f4",x"0e",x"5d",x"5c"),
   575 => (x"59",x"a6",x"cc",x"86"),
   576 => (x"c5",x"05",x"66",x"c8"),
   577 => (x"c3",x"48",x"c0",x"87"),
   578 => (x"66",x"c8",x"87",x"c7"),
   579 => (x"70",x"80",x"c8",x"48"),
   580 => (x"78",x"c0",x"48",x"7e"),
   581 => (x"c7",x"02",x"66",x"dc"),
   582 => (x"97",x"66",x"dc",x"87"),
   583 => (x"87",x"c5",x"05",x"bf"),
   584 => (x"ec",x"c2",x"48",x"c0"),
   585 => (x"c1",x"1e",x"c0",x"87"),
   586 => (x"e9",x"ca",x"49",x"49"),
   587 => (x"70",x"86",x"c4",x"87"),
   588 => (x"c0",x"02",x"9c",x"4c"),
   589 => (x"eb",x"c2",x"87",x"fc"),
   590 => (x"66",x"dc",x"4a",x"fc"),
   591 => (x"ca",x"de",x"ff",x"49"),
   592 => (x"02",x"98",x"70",x"87"),
   593 => (x"74",x"87",x"eb",x"c0"),
   594 => (x"49",x"66",x"dc",x"4a"),
   595 => (x"de",x"ff",x"4b",x"cb"),
   596 => (x"98",x"70",x"87",x"ee"),
   597 => (x"c0",x"87",x"db",x"02"),
   598 => (x"02",x"9c",x"74",x"1e"),
   599 => (x"4d",x"c0",x"87",x"c4"),
   600 => (x"4d",x"c1",x"87",x"c2"),
   601 => (x"ed",x"c9",x"49",x"75"),
   602 => (x"70",x"86",x"c4",x"87"),
   603 => (x"ff",x"05",x"9c",x"4c"),
   604 => (x"9c",x"74",x"87",x"c4"),
   605 => (x"87",x"d7",x"c1",x"02"),
   606 => (x"6e",x"49",x"a4",x"dc"),
   607 => (x"da",x"78",x"69",x"48"),
   608 => (x"66",x"c8",x"49",x"a4"),
   609 => (x"c8",x"80",x"c4",x"48"),
   610 => (x"69",x"9f",x"58",x"a6"),
   611 => (x"08",x"66",x"c4",x"48"),
   612 => (x"f4",x"eb",x"c2",x"78"),
   613 => (x"87",x"d2",x"02",x"bf"),
   614 => (x"9f",x"49",x"a4",x"d4"),
   615 => (x"ff",x"c0",x"49",x"69"),
   616 => (x"48",x"71",x"99",x"ff"),
   617 => (x"7e",x"70",x"30",x"d0"),
   618 => (x"7e",x"c0",x"87",x"c2"),
   619 => (x"66",x"c4",x"48",x"6e"),
   620 => (x"66",x"c4",x"80",x"bf"),
   621 => (x"66",x"c8",x"78",x"08"),
   622 => (x"c8",x"78",x"c0",x"48"),
   623 => (x"81",x"cc",x"49",x"66"),
   624 => (x"79",x"bf",x"66",x"c4"),
   625 => (x"d0",x"49",x"66",x"c8"),
   626 => (x"c1",x"79",x"c0",x"81"),
   627 => (x"c0",x"87",x"c2",x"48"),
   628 => (x"26",x"8e",x"f4",x"48"),
   629 => (x"26",x"4c",x"26",x"4d"),
   630 => (x"0e",x"4f",x"26",x"4b"),
   631 => (x"5d",x"5c",x"5b",x"5e"),
   632 => (x"d0",x"4c",x"71",x"0e"),
   633 => (x"9c",x"74",x"4d",x"66"),
   634 => (x"87",x"c2",x"c1",x"02"),
   635 => (x"69",x"49",x"a4",x"c8"),
   636 => (x"87",x"fa",x"c0",x"02"),
   637 => (x"75",x"85",x"49",x"6c"),
   638 => (x"f0",x"eb",x"c2",x"b9"),
   639 => (x"ba",x"ff",x"4a",x"bf"),
   640 => (x"99",x"71",x"99",x"72"),
   641 => (x"87",x"e4",x"c0",x"02"),
   642 => (x"6b",x"4b",x"a4",x"c4"),
   643 => (x"87",x"ee",x"f9",x"49"),
   644 => (x"eb",x"c2",x"7b",x"70"),
   645 => (x"6c",x"49",x"bf",x"ec"),
   646 => (x"75",x"7c",x"71",x"81"),
   647 => (x"f0",x"eb",x"c2",x"b9"),
   648 => (x"ba",x"ff",x"4a",x"bf"),
   649 => (x"99",x"71",x"99",x"72"),
   650 => (x"87",x"dc",x"ff",x"05"),
   651 => (x"4d",x"26",x"7c",x"75"),
   652 => (x"4b",x"26",x"4c",x"26"),
   653 => (x"73",x"1e",x"4f",x"26"),
   654 => (x"9b",x"4b",x"71",x"1e"),
   655 => (x"c8",x"87",x"c7",x"02"),
   656 => (x"05",x"69",x"49",x"a3"),
   657 => (x"48",x"c0",x"87",x"c5"),
   658 => (x"c2",x"87",x"f6",x"c0"),
   659 => (x"49",x"bf",x"c8",x"f0"),
   660 => (x"6a",x"4a",x"a3",x"c4"),
   661 => (x"c2",x"8a",x"c2",x"4a"),
   662 => (x"92",x"bf",x"ec",x"eb"),
   663 => (x"c2",x"49",x"a1",x"72"),
   664 => (x"4a",x"bf",x"f0",x"eb"),
   665 => (x"a1",x"72",x"9a",x"6b"),
   666 => (x"d4",x"f7",x"c0",x"49"),
   667 => (x"1e",x"66",x"c8",x"59"),
   668 => (x"87",x"cc",x"ea",x"71"),
   669 => (x"98",x"70",x"86",x"c4"),
   670 => (x"c0",x"87",x"c4",x"05"),
   671 => (x"c1",x"87",x"c2",x"48"),
   672 => (x"26",x"4b",x"26",x"48"),
   673 => (x"1e",x"73",x"1e",x"4f"),
   674 => (x"02",x"9b",x"4b",x"71"),
   675 => (x"a3",x"c8",x"87",x"c7"),
   676 => (x"c5",x"05",x"69",x"49"),
   677 => (x"c0",x"48",x"c0",x"87"),
   678 => (x"f0",x"c2",x"87",x"f6"),
   679 => (x"c4",x"49",x"bf",x"c8"),
   680 => (x"4a",x"6a",x"4a",x"a3"),
   681 => (x"eb",x"c2",x"8a",x"c2"),
   682 => (x"72",x"92",x"bf",x"ec"),
   683 => (x"eb",x"c2",x"49",x"a1"),
   684 => (x"6b",x"4a",x"bf",x"f0"),
   685 => (x"49",x"a1",x"72",x"9a"),
   686 => (x"59",x"d4",x"f7",x"c0"),
   687 => (x"71",x"1e",x"66",x"c8"),
   688 => (x"c4",x"87",x"d9",x"e5"),
   689 => (x"05",x"98",x"70",x"86"),
   690 => (x"48",x"c0",x"87",x"c4"),
   691 => (x"48",x"c1",x"87",x"c2"),
   692 => (x"4f",x"26",x"4b",x"26"),
   693 => (x"5c",x"5b",x"5e",x"0e"),
   694 => (x"86",x"fc",x"0e",x"5d"),
   695 => (x"66",x"d4",x"4b",x"71"),
   696 => (x"02",x"9b",x"73",x"4d"),
   697 => (x"c8",x"87",x"cc",x"c1"),
   698 => (x"02",x"69",x"49",x"a3"),
   699 => (x"d0",x"87",x"c4",x"c1"),
   700 => (x"eb",x"c2",x"4c",x"a3"),
   701 => (x"ff",x"49",x"bf",x"f0"),
   702 => (x"99",x"4a",x"6c",x"b9"),
   703 => (x"a9",x"66",x"d4",x"7e"),
   704 => (x"c0",x"87",x"cd",x"06"),
   705 => (x"a3",x"cc",x"7c",x"7b"),
   706 => (x"49",x"a3",x"c4",x"4a"),
   707 => (x"87",x"ca",x"79",x"6a"),
   708 => (x"c0",x"f8",x"49",x"72"),
   709 => (x"4d",x"66",x"d4",x"99"),
   710 => (x"49",x"75",x"8d",x"71"),
   711 => (x"1e",x"71",x"29",x"c9"),
   712 => (x"f6",x"fa",x"49",x"73"),
   713 => (x"ec",x"e3",x"c2",x"87"),
   714 => (x"fc",x"49",x"73",x"1e"),
   715 => (x"86",x"c8",x"87",x"c8"),
   716 => (x"fc",x"7c",x"66",x"d4"),
   717 => (x"26",x"4d",x"26",x"8e"),
   718 => (x"26",x"4b",x"26",x"4c"),
   719 => (x"1e",x"73",x"1e",x"4f"),
   720 => (x"02",x"9b",x"4b",x"71"),
   721 => (x"c2",x"87",x"e4",x"c0"),
   722 => (x"73",x"5b",x"dc",x"f0"),
   723 => (x"c2",x"8a",x"c2",x"4a"),
   724 => (x"49",x"bf",x"ec",x"eb"),
   725 => (x"c8",x"f0",x"c2",x"92"),
   726 => (x"80",x"72",x"48",x"bf"),
   727 => (x"58",x"e0",x"f0",x"c2"),
   728 => (x"30",x"c4",x"48",x"71"),
   729 => (x"58",x"fc",x"eb",x"c2"),
   730 => (x"c2",x"87",x"ed",x"c0"),
   731 => (x"c2",x"48",x"d8",x"f0"),
   732 => (x"78",x"bf",x"cc",x"f0"),
   733 => (x"48",x"dc",x"f0",x"c2"),
   734 => (x"bf",x"d0",x"f0",x"c2"),
   735 => (x"f4",x"eb",x"c2",x"78"),
   736 => (x"87",x"c9",x"02",x"bf"),
   737 => (x"bf",x"ec",x"eb",x"c2"),
   738 => (x"c7",x"31",x"c4",x"49"),
   739 => (x"d4",x"f0",x"c2",x"87"),
   740 => (x"31",x"c4",x"49",x"bf"),
   741 => (x"59",x"fc",x"eb",x"c2"),
   742 => (x"4f",x"26",x"4b",x"26"),
   743 => (x"5c",x"5b",x"5e",x"0e"),
   744 => (x"c0",x"4a",x"71",x"0e"),
   745 => (x"02",x"9a",x"72",x"4b"),
   746 => (x"da",x"87",x"e0",x"c0"),
   747 => (x"69",x"9f",x"49",x"a2"),
   748 => (x"f4",x"eb",x"c2",x"4b"),
   749 => (x"87",x"cf",x"02",x"bf"),
   750 => (x"9f",x"49",x"a2",x"d4"),
   751 => (x"c0",x"4c",x"49",x"69"),
   752 => (x"d0",x"9c",x"ff",x"ff"),
   753 => (x"c0",x"87",x"c2",x"34"),
   754 => (x"73",x"b3",x"74",x"4c"),
   755 => (x"87",x"ed",x"fd",x"49"),
   756 => (x"4b",x"26",x"4c",x"26"),
   757 => (x"5e",x"0e",x"4f",x"26"),
   758 => (x"0e",x"5d",x"5c",x"5b"),
   759 => (x"a6",x"c8",x"86",x"f0"),
   760 => (x"ff",x"ff",x"cf",x"59"),
   761 => (x"c0",x"4c",x"f8",x"ff"),
   762 => (x"02",x"66",x"c4",x"7e"),
   763 => (x"e3",x"c2",x"87",x"d8"),
   764 => (x"78",x"c0",x"48",x"e8"),
   765 => (x"48",x"e0",x"e3",x"c2"),
   766 => (x"bf",x"dc",x"f0",x"c2"),
   767 => (x"e4",x"e3",x"c2",x"78"),
   768 => (x"d8",x"f0",x"c2",x"48"),
   769 => (x"ec",x"c2",x"78",x"bf"),
   770 => (x"50",x"c0",x"48",x"c9"),
   771 => (x"bf",x"f8",x"eb",x"c2"),
   772 => (x"e8",x"e3",x"c2",x"49"),
   773 => (x"aa",x"71",x"4a",x"bf"),
   774 => (x"87",x"cb",x"c4",x"03"),
   775 => (x"99",x"cf",x"49",x"72"),
   776 => (x"87",x"e9",x"c0",x"05"),
   777 => (x"48",x"d0",x"f7",x"c0"),
   778 => (x"bf",x"e0",x"e3",x"c2"),
   779 => (x"ec",x"e3",x"c2",x"78"),
   780 => (x"e0",x"e3",x"c2",x"1e"),
   781 => (x"e3",x"c2",x"49",x"bf"),
   782 => (x"a1",x"c1",x"48",x"e0"),
   783 => (x"ff",x"e2",x"71",x"78"),
   784 => (x"c0",x"86",x"c4",x"87"),
   785 => (x"c2",x"48",x"cc",x"f7"),
   786 => (x"cc",x"78",x"ec",x"e3"),
   787 => (x"cc",x"f7",x"c0",x"87"),
   788 => (x"e0",x"c0",x"48",x"bf"),
   789 => (x"d0",x"f7",x"c0",x"80"),
   790 => (x"e8",x"e3",x"c2",x"58"),
   791 => (x"80",x"c1",x"48",x"bf"),
   792 => (x"58",x"ec",x"e3",x"c2"),
   793 => (x"00",x"0d",x"cc",x"27"),
   794 => (x"bf",x"97",x"bf",x"00"),
   795 => (x"c2",x"02",x"9d",x"4d"),
   796 => (x"e5",x"c3",x"87",x"e5"),
   797 => (x"de",x"c2",x"02",x"ad"),
   798 => (x"cc",x"f7",x"c0",x"87"),
   799 => (x"a3",x"cb",x"4b",x"bf"),
   800 => (x"cf",x"4c",x"11",x"49"),
   801 => (x"d2",x"c1",x"05",x"ac"),
   802 => (x"df",x"49",x"75",x"87"),
   803 => (x"cd",x"89",x"c1",x"99"),
   804 => (x"fc",x"eb",x"c2",x"91"),
   805 => (x"4a",x"a3",x"c1",x"81"),
   806 => (x"a3",x"c3",x"51",x"12"),
   807 => (x"c5",x"51",x"12",x"4a"),
   808 => (x"51",x"12",x"4a",x"a3"),
   809 => (x"12",x"4a",x"a3",x"c7"),
   810 => (x"4a",x"a3",x"c9",x"51"),
   811 => (x"a3",x"ce",x"51",x"12"),
   812 => (x"d0",x"51",x"12",x"4a"),
   813 => (x"51",x"12",x"4a",x"a3"),
   814 => (x"12",x"4a",x"a3",x"d2"),
   815 => (x"4a",x"a3",x"d4",x"51"),
   816 => (x"a3",x"d6",x"51",x"12"),
   817 => (x"d8",x"51",x"12",x"4a"),
   818 => (x"51",x"12",x"4a",x"a3"),
   819 => (x"12",x"4a",x"a3",x"dc"),
   820 => (x"4a",x"a3",x"de",x"51"),
   821 => (x"7e",x"c1",x"51",x"12"),
   822 => (x"74",x"87",x"fc",x"c0"),
   823 => (x"05",x"99",x"c8",x"49"),
   824 => (x"74",x"87",x"ed",x"c0"),
   825 => (x"05",x"99",x"d0",x"49"),
   826 => (x"e0",x"c0",x"87",x"d3"),
   827 => (x"cc",x"c0",x"02",x"66"),
   828 => (x"c0",x"49",x"73",x"87"),
   829 => (x"70",x"0f",x"66",x"e0"),
   830 => (x"d3",x"c0",x"02",x"98"),
   831 => (x"c0",x"05",x"6e",x"87"),
   832 => (x"eb",x"c2",x"87",x"c6"),
   833 => (x"50",x"c0",x"48",x"fc"),
   834 => (x"bf",x"cc",x"f7",x"c0"),
   835 => (x"87",x"e9",x"c2",x"48"),
   836 => (x"48",x"c9",x"ec",x"c2"),
   837 => (x"c2",x"7e",x"50",x"c0"),
   838 => (x"49",x"bf",x"f8",x"eb"),
   839 => (x"bf",x"e8",x"e3",x"c2"),
   840 => (x"04",x"aa",x"71",x"4a"),
   841 => (x"cf",x"87",x"f5",x"fb"),
   842 => (x"f8",x"ff",x"ff",x"ff"),
   843 => (x"dc",x"f0",x"c2",x"4c"),
   844 => (x"c8",x"c0",x"05",x"bf"),
   845 => (x"f4",x"eb",x"c2",x"87"),
   846 => (x"fa",x"c1",x"02",x"bf"),
   847 => (x"e4",x"e3",x"c2",x"87"),
   848 => (x"f9",x"ec",x"49",x"bf"),
   849 => (x"e8",x"e3",x"c2",x"87"),
   850 => (x"48",x"a6",x"c4",x"58"),
   851 => (x"bf",x"e4",x"e3",x"c2"),
   852 => (x"f4",x"eb",x"c2",x"78"),
   853 => (x"db",x"c0",x"02",x"bf"),
   854 => (x"49",x"66",x"c4",x"87"),
   855 => (x"a9",x"74",x"99",x"74"),
   856 => (x"87",x"c8",x"c0",x"02"),
   857 => (x"c0",x"48",x"a6",x"c8"),
   858 => (x"87",x"e7",x"c0",x"78"),
   859 => (x"c1",x"48",x"a6",x"c8"),
   860 => (x"87",x"df",x"c0",x"78"),
   861 => (x"cf",x"49",x"66",x"c4"),
   862 => (x"a9",x"99",x"f8",x"ff"),
   863 => (x"87",x"c8",x"c0",x"02"),
   864 => (x"c0",x"48",x"a6",x"cc"),
   865 => (x"87",x"c5",x"c0",x"78"),
   866 => (x"c1",x"48",x"a6",x"cc"),
   867 => (x"48",x"a6",x"c8",x"78"),
   868 => (x"c8",x"78",x"66",x"cc"),
   869 => (x"de",x"c0",x"05",x"66"),
   870 => (x"49",x"66",x"c4",x"87"),
   871 => (x"eb",x"c2",x"89",x"c2"),
   872 => (x"c2",x"91",x"bf",x"ec"),
   873 => (x"48",x"bf",x"c8",x"f0"),
   874 => (x"e3",x"c2",x"80",x"71"),
   875 => (x"e3",x"c2",x"58",x"e4"),
   876 => (x"78",x"c0",x"48",x"e8"),
   877 => (x"c0",x"87",x"d5",x"f9"),
   878 => (x"ff",x"ff",x"cf",x"48"),
   879 => (x"f0",x"4c",x"f8",x"ff"),
   880 => (x"26",x"4d",x"26",x"8e"),
   881 => (x"26",x"4b",x"26",x"4c"),
   882 => (x"00",x"00",x"00",x"4f"),
   883 => (x"00",x"00",x"00",x"00"),
   884 => (x"ff",x"ff",x"ff",x"ff"),
   885 => (x"00",x"00",x"0d",x"dc"),
   886 => (x"00",x"00",x"0d",x"e8"),
   887 => (x"33",x"54",x"41",x"46"),
   888 => (x"20",x"20",x"20",x"32"),
   889 => (x"00",x"00",x"00",x"00"),
   890 => (x"31",x"54",x"41",x"46"),
   891 => (x"20",x"20",x"20",x"36"),
   892 => (x"d4",x"ff",x"1e",x"00"),
   893 => (x"78",x"ff",x"c3",x"48"),
   894 => (x"4f",x"26",x"48",x"68"),
   895 => (x"48",x"d4",x"ff",x"1e"),
   896 => (x"ff",x"78",x"ff",x"c3"),
   897 => (x"e1",x"c0",x"48",x"d0"),
   898 => (x"48",x"d4",x"ff",x"78"),
   899 => (x"4f",x"26",x"78",x"d4"),
   900 => (x"48",x"d0",x"ff",x"1e"),
   901 => (x"26",x"78",x"e0",x"c0"),
   902 => (x"d4",x"ff",x"1e",x"4f"),
   903 => (x"99",x"49",x"70",x"87"),
   904 => (x"c0",x"87",x"c6",x"02"),
   905 => (x"f1",x"05",x"a9",x"fb"),
   906 => (x"26",x"48",x"71",x"87"),
   907 => (x"5b",x"5e",x"0e",x"4f"),
   908 => (x"4b",x"71",x"0e",x"5c"),
   909 => (x"f8",x"fe",x"4c",x"c0"),
   910 => (x"99",x"49",x"70",x"87"),
   911 => (x"87",x"f9",x"c0",x"02"),
   912 => (x"02",x"a9",x"ec",x"c0"),
   913 => (x"c0",x"87",x"f2",x"c0"),
   914 => (x"c0",x"02",x"a9",x"fb"),
   915 => (x"66",x"cc",x"87",x"eb"),
   916 => (x"c7",x"03",x"ac",x"b7"),
   917 => (x"02",x"66",x"d0",x"87"),
   918 => (x"53",x"71",x"87",x"c2"),
   919 => (x"c2",x"02",x"99",x"71"),
   920 => (x"fe",x"84",x"c1",x"87"),
   921 => (x"49",x"70",x"87",x"cb"),
   922 => (x"87",x"cd",x"02",x"99"),
   923 => (x"02",x"a9",x"ec",x"c0"),
   924 => (x"fb",x"c0",x"87",x"c7"),
   925 => (x"d5",x"ff",x"05",x"a9"),
   926 => (x"02",x"66",x"d0",x"87"),
   927 => (x"97",x"c0",x"87",x"c3"),
   928 => (x"a9",x"ec",x"c0",x"7b"),
   929 => (x"74",x"87",x"c4",x"05"),
   930 => (x"74",x"87",x"c5",x"4a"),
   931 => (x"8a",x"0a",x"c0",x"4a"),
   932 => (x"4c",x"26",x"48",x"72"),
   933 => (x"4f",x"26",x"4b",x"26"),
   934 => (x"87",x"d5",x"fd",x"1e"),
   935 => (x"f0",x"c0",x"49",x"70"),
   936 => (x"87",x"c9",x"04",x"a9"),
   937 => (x"01",x"a9",x"f9",x"c0"),
   938 => (x"f0",x"c0",x"87",x"c3"),
   939 => (x"a9",x"c1",x"c1",x"89"),
   940 => (x"c1",x"87",x"c9",x"04"),
   941 => (x"c3",x"01",x"a9",x"da"),
   942 => (x"89",x"f7",x"c0",x"87"),
   943 => (x"4f",x"26",x"48",x"71"),
   944 => (x"5c",x"5b",x"5e",x"0e"),
   945 => (x"86",x"f8",x"0e",x"5d"),
   946 => (x"7e",x"c0",x"4c",x"71"),
   947 => (x"c0",x"87",x"ed",x"fc"),
   948 => (x"e0",x"fd",x"c0",x"4b"),
   949 => (x"c0",x"49",x"bf",x"97"),
   950 => (x"87",x"cf",x"04",x"a9"),
   951 => (x"c1",x"87",x"fa",x"fc"),
   952 => (x"e0",x"fd",x"c0",x"83"),
   953 => (x"ab",x"49",x"bf",x"97"),
   954 => (x"c0",x"87",x"f1",x"06"),
   955 => (x"bf",x"97",x"e0",x"fd"),
   956 => (x"fb",x"87",x"cf",x"02"),
   957 => (x"49",x"70",x"87",x"fb"),
   958 => (x"87",x"c6",x"02",x"99"),
   959 => (x"05",x"a9",x"ec",x"c0"),
   960 => (x"4b",x"c0",x"87",x"f1"),
   961 => (x"70",x"87",x"ea",x"fb"),
   962 => (x"87",x"e5",x"fb",x"4d"),
   963 => (x"fb",x"58",x"a6",x"c8"),
   964 => (x"4a",x"70",x"87",x"df"),
   965 => (x"a4",x"c8",x"83",x"c1"),
   966 => (x"49",x"69",x"97",x"49"),
   967 => (x"87",x"da",x"05",x"ad"),
   968 => (x"97",x"49",x"a4",x"c9"),
   969 => (x"66",x"c4",x"49",x"69"),
   970 => (x"87",x"ce",x"05",x"a9"),
   971 => (x"97",x"49",x"a4",x"ca"),
   972 => (x"05",x"aa",x"49",x"69"),
   973 => (x"7e",x"c1",x"87",x"c4"),
   974 => (x"ec",x"c0",x"87",x"d0"),
   975 => (x"87",x"c6",x"02",x"ad"),
   976 => (x"05",x"ad",x"fb",x"c0"),
   977 => (x"4b",x"c0",x"87",x"c4"),
   978 => (x"02",x"6e",x"7e",x"c1"),
   979 => (x"fa",x"87",x"f5",x"fe"),
   980 => (x"48",x"73",x"87",x"fe"),
   981 => (x"4d",x"26",x"8e",x"f8"),
   982 => (x"4b",x"26",x"4c",x"26"),
   983 => (x"00",x"00",x"4f",x"26"),
   984 => (x"1e",x"73",x"1e",x"00"),
   985 => (x"c8",x"4b",x"d4",x"ff"),
   986 => (x"d0",x"ff",x"4a",x"66"),
   987 => (x"78",x"c5",x"c8",x"48"),
   988 => (x"c1",x"48",x"d4",x"ff"),
   989 => (x"7b",x"11",x"78",x"d4"),
   990 => (x"f9",x"05",x"8a",x"c1"),
   991 => (x"48",x"d0",x"ff",x"87"),
   992 => (x"4b",x"26",x"78",x"c4"),
   993 => (x"5e",x"0e",x"4f",x"26"),
   994 => (x"0e",x"5d",x"5c",x"5b"),
   995 => (x"7e",x"71",x"86",x"f8"),
   996 => (x"f0",x"c2",x"1e",x"6e"),
   997 => (x"dc",x"e5",x"49",x"ec"),
   998 => (x"70",x"86",x"c4",x"87"),
   999 => (x"e4",x"c4",x"02",x"98"),
  1000 => (x"e8",x"ec",x"c1",x"87"),
  1001 => (x"49",x"6e",x"4c",x"bf"),
  1002 => (x"c8",x"87",x"d5",x"fc"),
  1003 => (x"98",x"70",x"58",x"a6"),
  1004 => (x"c4",x"87",x"c5",x"05"),
  1005 => (x"78",x"c1",x"48",x"a6"),
  1006 => (x"c5",x"48",x"d0",x"ff"),
  1007 => (x"48",x"d4",x"ff",x"78"),
  1008 => (x"c4",x"78",x"d5",x"c1"),
  1009 => (x"89",x"c1",x"49",x"66"),
  1010 => (x"ec",x"c1",x"31",x"c6"),
  1011 => (x"4a",x"bf",x"97",x"e0"),
  1012 => (x"ff",x"b0",x"71",x"48"),
  1013 => (x"ff",x"78",x"08",x"d4"),
  1014 => (x"78",x"c4",x"48",x"d0"),
  1015 => (x"97",x"e8",x"f0",x"c2"),
  1016 => (x"99",x"d0",x"49",x"bf"),
  1017 => (x"c5",x"87",x"dd",x"02"),
  1018 => (x"48",x"d4",x"ff",x"78"),
  1019 => (x"c0",x"78",x"d6",x"c1"),
  1020 => (x"48",x"d4",x"ff",x"4a"),
  1021 => (x"c1",x"78",x"ff",x"c3"),
  1022 => (x"aa",x"e0",x"c0",x"82"),
  1023 => (x"ff",x"87",x"f2",x"04"),
  1024 => (x"78",x"c4",x"48",x"d0"),
  1025 => (x"c3",x"48",x"d4",x"ff"),
  1026 => (x"d0",x"ff",x"78",x"ff"),
  1027 => (x"ff",x"78",x"c5",x"48"),
  1028 => (x"d3",x"c1",x"48",x"d4"),
  1029 => (x"ff",x"78",x"c1",x"78"),
  1030 => (x"78",x"c4",x"48",x"d0"),
  1031 => (x"06",x"ac",x"b7",x"c0"),
  1032 => (x"c2",x"87",x"cb",x"c2"),
  1033 => (x"4b",x"bf",x"f4",x"f0"),
  1034 => (x"73",x"7e",x"74",x"8c"),
  1035 => (x"dd",x"c1",x"02",x"9b"),
  1036 => (x"4d",x"c0",x"c8",x"87"),
  1037 => (x"ab",x"b7",x"c0",x"8b"),
  1038 => (x"c8",x"87",x"c6",x"03"),
  1039 => (x"c0",x"4d",x"a3",x"c0"),
  1040 => (x"e8",x"f0",x"c2",x"4b"),
  1041 => (x"d0",x"49",x"bf",x"97"),
  1042 => (x"87",x"cf",x"02",x"99"),
  1043 => (x"f0",x"c2",x"1e",x"c0"),
  1044 => (x"e1",x"e7",x"49",x"ec"),
  1045 => (x"70",x"86",x"c4",x"87"),
  1046 => (x"c2",x"87",x"d8",x"4c"),
  1047 => (x"c2",x"1e",x"ec",x"e3"),
  1048 => (x"e7",x"49",x"ec",x"f0"),
  1049 => (x"4c",x"70",x"87",x"d0"),
  1050 => (x"e3",x"c2",x"1e",x"75"),
  1051 => (x"f0",x"fb",x"49",x"ec"),
  1052 => (x"74",x"86",x"c8",x"87"),
  1053 => (x"87",x"c5",x"05",x"9c"),
  1054 => (x"ca",x"c1",x"48",x"c0"),
  1055 => (x"c2",x"1e",x"c1",x"87"),
  1056 => (x"e5",x"49",x"ec",x"f0"),
  1057 => (x"86",x"c4",x"87",x"d5"),
  1058 => (x"fe",x"05",x"9b",x"73"),
  1059 => (x"4c",x"6e",x"87",x"e3"),
  1060 => (x"06",x"ac",x"b7",x"c0"),
  1061 => (x"f0",x"c2",x"87",x"d1"),
  1062 => (x"78",x"c0",x"48",x"ec"),
  1063 => (x"78",x"c0",x"80",x"d0"),
  1064 => (x"f0",x"c2",x"80",x"f4"),
  1065 => (x"c0",x"78",x"bf",x"f8"),
  1066 => (x"fd",x"01",x"ac",x"b7"),
  1067 => (x"d0",x"ff",x"87",x"f5"),
  1068 => (x"ff",x"78",x"c5",x"48"),
  1069 => (x"d3",x"c1",x"48",x"d4"),
  1070 => (x"ff",x"78",x"c0",x"78"),
  1071 => (x"78",x"c4",x"48",x"d0"),
  1072 => (x"c2",x"c0",x"48",x"c1"),
  1073 => (x"f8",x"48",x"c0",x"87"),
  1074 => (x"26",x"4d",x"26",x"8e"),
  1075 => (x"26",x"4b",x"26",x"4c"),
  1076 => (x"5b",x"5e",x"0e",x"4f"),
  1077 => (x"fc",x"0e",x"5d",x"5c"),
  1078 => (x"c0",x"4d",x"71",x"86"),
  1079 => (x"04",x"ad",x"4c",x"4b"),
  1080 => (x"c0",x"87",x"e8",x"c0"),
  1081 => (x"74",x"1e",x"c0",x"fb"),
  1082 => (x"87",x"c4",x"02",x"9c"),
  1083 => (x"87",x"c2",x"4a",x"c0"),
  1084 => (x"49",x"72",x"4a",x"c1"),
  1085 => (x"c4",x"87",x"df",x"eb"),
  1086 => (x"c1",x"7e",x"70",x"86"),
  1087 => (x"c2",x"05",x"6e",x"83"),
  1088 => (x"c1",x"4b",x"75",x"87"),
  1089 => (x"06",x"ab",x"75",x"84"),
  1090 => (x"6e",x"87",x"d8",x"ff"),
  1091 => (x"26",x"8e",x"fc",x"48"),
  1092 => (x"26",x"4c",x"26",x"4d"),
  1093 => (x"0e",x"4f",x"26",x"4b"),
  1094 => (x"0e",x"5c",x"5b",x"5e"),
  1095 => (x"66",x"cc",x"4b",x"71"),
  1096 => (x"4c",x"87",x"d8",x"02"),
  1097 => (x"02",x"8c",x"f0",x"c0"),
  1098 => (x"4a",x"74",x"87",x"d8"),
  1099 => (x"d1",x"02",x"8a",x"c1"),
  1100 => (x"cd",x"02",x"8a",x"87"),
  1101 => (x"c9",x"02",x"8a",x"87"),
  1102 => (x"73",x"87",x"d9",x"87"),
  1103 => (x"87",x"c6",x"f9",x"49"),
  1104 => (x"1e",x"74",x"87",x"d2"),
  1105 => (x"da",x"c1",x"49",x"c0"),
  1106 => (x"1e",x"74",x"87",x"e2"),
  1107 => (x"da",x"c1",x"49",x"73"),
  1108 => (x"86",x"c8",x"87",x"da"),
  1109 => (x"4b",x"26",x"4c",x"26"),
  1110 => (x"5e",x"0e",x"4f",x"26"),
  1111 => (x"0e",x"5d",x"5c",x"5b"),
  1112 => (x"4c",x"71",x"86",x"fc"),
  1113 => (x"c2",x"91",x"de",x"49"),
  1114 => (x"71",x"4d",x"d8",x"f1"),
  1115 => (x"02",x"6d",x"97",x"85"),
  1116 => (x"c2",x"87",x"dc",x"c1"),
  1117 => (x"49",x"bf",x"c8",x"f1"),
  1118 => (x"fd",x"71",x"81",x"74"),
  1119 => (x"7e",x"70",x"87",x"d3"),
  1120 => (x"c0",x"02",x"98",x"48"),
  1121 => (x"f1",x"c2",x"87",x"f2"),
  1122 => (x"4a",x"70",x"4b",x"cc"),
  1123 => (x"fe",x"fe",x"49",x"cb"),
  1124 => (x"4b",x"74",x"87",x"d2"),
  1125 => (x"ec",x"c1",x"93",x"cc"),
  1126 => (x"83",x"c4",x"83",x"ec"),
  1127 => (x"7b",x"dc",x"c7",x"c1"),
  1128 => (x"c4",x"c1",x"49",x"74"),
  1129 => (x"7b",x"75",x"87",x"da"),
  1130 => (x"97",x"e4",x"ec",x"c1"),
  1131 => (x"c2",x"1e",x"49",x"bf"),
  1132 => (x"fd",x"49",x"cc",x"f1"),
  1133 => (x"86",x"c4",x"87",x"e1"),
  1134 => (x"c4",x"c1",x"49",x"74"),
  1135 => (x"49",x"c0",x"87",x"c2"),
  1136 => (x"87",x"dd",x"c5",x"c1"),
  1137 => (x"48",x"e4",x"f0",x"c2"),
  1138 => (x"c0",x"49",x"50",x"c0"),
  1139 => (x"fc",x"87",x"cc",x"e2"),
  1140 => (x"26",x"4d",x"26",x"8e"),
  1141 => (x"26",x"4b",x"26",x"4c"),
  1142 => (x"00",x"00",x"00",x"4f"),
  1143 => (x"64",x"61",x"6f",x"4c"),
  1144 => (x"2e",x"67",x"6e",x"69"),
  1145 => (x"1e",x"00",x"2e",x"2e"),
  1146 => (x"4b",x"71",x"1e",x"73"),
  1147 => (x"c8",x"f1",x"c2",x"49"),
  1148 => (x"fb",x"71",x"81",x"bf"),
  1149 => (x"4a",x"70",x"87",x"db"),
  1150 => (x"87",x"c4",x"02",x"9a"),
  1151 => (x"87",x"dc",x"e6",x"49"),
  1152 => (x"48",x"c8",x"f1",x"c2"),
  1153 => (x"49",x"73",x"78",x"c0"),
  1154 => (x"26",x"87",x"fa",x"c1"),
  1155 => (x"1e",x"4f",x"26",x"4b"),
  1156 => (x"4b",x"71",x"1e",x"73"),
  1157 => (x"02",x"4a",x"a3",x"c4"),
  1158 => (x"c1",x"87",x"d0",x"c1"),
  1159 => (x"87",x"dc",x"02",x"8a"),
  1160 => (x"f2",x"c0",x"02",x"8a"),
  1161 => (x"c1",x"05",x"8a",x"87"),
  1162 => (x"f1",x"c2",x"87",x"d3"),
  1163 => (x"c1",x"02",x"bf",x"c8"),
  1164 => (x"c1",x"48",x"87",x"cb"),
  1165 => (x"cc",x"f1",x"c2",x"88"),
  1166 => (x"87",x"c1",x"c1",x"58"),
  1167 => (x"bf",x"c8",x"f1",x"c2"),
  1168 => (x"c2",x"89",x"c6",x"49"),
  1169 => (x"c0",x"59",x"cc",x"f1"),
  1170 => (x"c0",x"03",x"a9",x"b7"),
  1171 => (x"f1",x"c2",x"87",x"ef"),
  1172 => (x"78",x"c0",x"48",x"c8"),
  1173 => (x"c2",x"87",x"e6",x"c0"),
  1174 => (x"02",x"bf",x"c4",x"f1"),
  1175 => (x"f1",x"c2",x"87",x"df"),
  1176 => (x"c1",x"48",x"bf",x"c8"),
  1177 => (x"cc",x"f1",x"c2",x"80"),
  1178 => (x"c2",x"87",x"d2",x"58"),
  1179 => (x"02",x"bf",x"c4",x"f1"),
  1180 => (x"f1",x"c2",x"87",x"cb"),
  1181 => (x"c6",x"48",x"bf",x"c8"),
  1182 => (x"cc",x"f1",x"c2",x"80"),
  1183 => (x"c4",x"49",x"73",x"58"),
  1184 => (x"26",x"4b",x"26",x"87"),
  1185 => (x"5b",x"5e",x"0e",x"4f"),
  1186 => (x"f0",x"0e",x"5d",x"5c"),
  1187 => (x"59",x"a6",x"d0",x"86"),
  1188 => (x"4d",x"ec",x"e3",x"c2"),
  1189 => (x"f1",x"c2",x"4c",x"c0"),
  1190 => (x"78",x"c1",x"48",x"c4"),
  1191 => (x"c0",x"48",x"a6",x"c8"),
  1192 => (x"c2",x"7e",x"75",x"78"),
  1193 => (x"48",x"bf",x"c8",x"f1"),
  1194 => (x"c1",x"06",x"a8",x"c0"),
  1195 => (x"a6",x"c8",x"87",x"c0"),
  1196 => (x"c2",x"7e",x"75",x"5c"),
  1197 => (x"98",x"48",x"ec",x"e3"),
  1198 => (x"87",x"f2",x"c0",x"02"),
  1199 => (x"c0",x"4d",x"66",x"c4"),
  1200 => (x"cc",x"1e",x"c0",x"fb"),
  1201 => (x"87",x"c4",x"02",x"66"),
  1202 => (x"87",x"c2",x"4c",x"c0"),
  1203 => (x"49",x"74",x"4c",x"c1"),
  1204 => (x"c4",x"87",x"c3",x"e4"),
  1205 => (x"c1",x"7e",x"70",x"86"),
  1206 => (x"48",x"66",x"c8",x"85"),
  1207 => (x"a6",x"cc",x"80",x"c1"),
  1208 => (x"c8",x"f1",x"c2",x"58"),
  1209 => (x"c5",x"03",x"ad",x"bf"),
  1210 => (x"ff",x"05",x"6e",x"87"),
  1211 => (x"4d",x"6e",x"87",x"d1"),
  1212 => (x"9d",x"75",x"4c",x"c0"),
  1213 => (x"87",x"dc",x"c3",x"02"),
  1214 => (x"1e",x"c0",x"fb",x"c0"),
  1215 => (x"c7",x"02",x"66",x"cc"),
  1216 => (x"48",x"a6",x"c8",x"87"),
  1217 => (x"87",x"c5",x"78",x"c0"),
  1218 => (x"c1",x"48",x"a6",x"c8"),
  1219 => (x"49",x"66",x"c8",x"78"),
  1220 => (x"c4",x"87",x"c3",x"e3"),
  1221 => (x"48",x"7e",x"70",x"86"),
  1222 => (x"e4",x"c2",x"02",x"98"),
  1223 => (x"81",x"cb",x"49",x"87"),
  1224 => (x"d0",x"49",x"69",x"97"),
  1225 => (x"d4",x"c1",x"02",x"99"),
  1226 => (x"cc",x"49",x"74",x"87"),
  1227 => (x"ec",x"ec",x"c1",x"91"),
  1228 => (x"e7",x"c7",x"c1",x"81"),
  1229 => (x"c3",x"81",x"c8",x"79"),
  1230 => (x"49",x"74",x"51",x"ff"),
  1231 => (x"f1",x"c2",x"91",x"de"),
  1232 => (x"85",x"71",x"4d",x"d8"),
  1233 => (x"7d",x"97",x"c1",x"c2"),
  1234 => (x"c0",x"49",x"a5",x"c1"),
  1235 => (x"eb",x"c2",x"51",x"e0"),
  1236 => (x"02",x"bf",x"97",x"fc"),
  1237 => (x"84",x"c1",x"87",x"d2"),
  1238 => (x"c2",x"4b",x"a5",x"c2"),
  1239 => (x"db",x"4a",x"fc",x"eb"),
  1240 => (x"ff",x"f6",x"fe",x"49"),
  1241 => (x"87",x"d9",x"c1",x"87"),
  1242 => (x"c0",x"49",x"a5",x"cd"),
  1243 => (x"c2",x"84",x"c1",x"51"),
  1244 => (x"4a",x"6e",x"4b",x"a5"),
  1245 => (x"f6",x"fe",x"49",x"cb"),
  1246 => (x"c4",x"c1",x"87",x"ea"),
  1247 => (x"cc",x"49",x"74",x"87"),
  1248 => (x"ec",x"ec",x"c1",x"91"),
  1249 => (x"da",x"c5",x"c1",x"81"),
  1250 => (x"fc",x"eb",x"c2",x"79"),
  1251 => (x"d8",x"02",x"bf",x"97"),
  1252 => (x"de",x"49",x"74",x"87"),
  1253 => (x"c2",x"84",x"c1",x"91"),
  1254 => (x"71",x"4b",x"d8",x"f1"),
  1255 => (x"fc",x"eb",x"c2",x"83"),
  1256 => (x"fe",x"49",x"dd",x"4a"),
  1257 => (x"d8",x"87",x"fd",x"f5"),
  1258 => (x"de",x"4b",x"74",x"87"),
  1259 => (x"d8",x"f1",x"c2",x"93"),
  1260 => (x"49",x"a3",x"cb",x"83"),
  1261 => (x"84",x"c1",x"51",x"c0"),
  1262 => (x"cb",x"4a",x"6e",x"73"),
  1263 => (x"e3",x"f5",x"fe",x"49"),
  1264 => (x"48",x"66",x"c8",x"87"),
  1265 => (x"a6",x"cc",x"80",x"c1"),
  1266 => (x"03",x"ac",x"c7",x"58"),
  1267 => (x"6e",x"87",x"c5",x"c0"),
  1268 => (x"87",x"e4",x"fc",x"05"),
  1269 => (x"c0",x"03",x"ac",x"c7"),
  1270 => (x"f1",x"c2",x"87",x"e4"),
  1271 => (x"78",x"c0",x"48",x"c4"),
  1272 => (x"91",x"cc",x"49",x"74"),
  1273 => (x"81",x"ec",x"ec",x"c1"),
  1274 => (x"79",x"da",x"c5",x"c1"),
  1275 => (x"91",x"de",x"49",x"74"),
  1276 => (x"81",x"d8",x"f1",x"c2"),
  1277 => (x"84",x"c1",x"51",x"c0"),
  1278 => (x"ff",x"04",x"ac",x"c7"),
  1279 => (x"ee",x"c1",x"87",x"dc"),
  1280 => (x"50",x"c0",x"48",x"c8"),
  1281 => (x"d1",x"c1",x"80",x"f7"),
  1282 => (x"d0",x"c1",x"40",x"f5"),
  1283 => (x"80",x"c8",x"78",x"e8"),
  1284 => (x"78",x"cf",x"c8",x"c1"),
  1285 => (x"c0",x"49",x"66",x"cc"),
  1286 => (x"f0",x"87",x"e5",x"fa"),
  1287 => (x"26",x"4d",x"26",x"8e"),
  1288 => (x"26",x"4b",x"26",x"4c"),
  1289 => (x"00",x"00",x"00",x"4f"),
  1290 => (x"61",x"42",x"20",x"80"),
  1291 => (x"1e",x"00",x"6b",x"63"),
  1292 => (x"4b",x"71",x"1e",x"73"),
  1293 => (x"c1",x"91",x"cc",x"49"),
  1294 => (x"c8",x"81",x"ec",x"ec"),
  1295 => (x"ec",x"c1",x"4a",x"a1"),
  1296 => (x"50",x"12",x"48",x"e0"),
  1297 => (x"c0",x"4a",x"a1",x"c9"),
  1298 => (x"12",x"48",x"e0",x"fd"),
  1299 => (x"c1",x"81",x"ca",x"50"),
  1300 => (x"11",x"48",x"e4",x"ec"),
  1301 => (x"e4",x"ec",x"c1",x"50"),
  1302 => (x"1e",x"49",x"bf",x"97"),
  1303 => (x"f6",x"f2",x"49",x"c0"),
  1304 => (x"f8",x"49",x"73",x"87"),
  1305 => (x"8e",x"fc",x"87",x"df"),
  1306 => (x"4f",x"26",x"4b",x"26"),
  1307 => (x"c0",x"49",x"c0",x"1e"),
  1308 => (x"26",x"87",x"ee",x"fa"),
  1309 => (x"4a",x"71",x"1e",x"4f"),
  1310 => (x"c1",x"91",x"cc",x"49"),
  1311 => (x"c8",x"81",x"ec",x"ec"),
  1312 => (x"e4",x"f0",x"c2",x"81"),
  1313 => (x"c0",x"50",x"11",x"48"),
  1314 => (x"fe",x"49",x"a2",x"f0"),
  1315 => (x"c0",x"87",x"fd",x"ef"),
  1316 => (x"87",x"c7",x"d7",x"49"),
  1317 => (x"ff",x"1e",x"4f",x"26"),
  1318 => (x"ff",x"c3",x"4a",x"d4"),
  1319 => (x"48",x"d0",x"ff",x"7a"),
  1320 => (x"de",x"78",x"e1",x"c0"),
  1321 => (x"48",x"7a",x"71",x"7a"),
  1322 => (x"70",x"28",x"b7",x"c8"),
  1323 => (x"d0",x"48",x"71",x"7a"),
  1324 => (x"7a",x"70",x"28",x"b7"),
  1325 => (x"b7",x"d8",x"48",x"71"),
  1326 => (x"ff",x"7a",x"70",x"28"),
  1327 => (x"e0",x"c0",x"48",x"d0"),
  1328 => (x"0e",x"4f",x"26",x"78"),
  1329 => (x"5d",x"5c",x"5b",x"5e"),
  1330 => (x"71",x"86",x"f4",x"0e"),
  1331 => (x"91",x"cc",x"49",x"4d"),
  1332 => (x"81",x"ec",x"ec",x"c1"),
  1333 => (x"ca",x"4a",x"a1",x"c8"),
  1334 => (x"a6",x"c4",x"7e",x"a1"),
  1335 => (x"e0",x"f0",x"c2",x"48"),
  1336 => (x"97",x"6e",x"78",x"bf"),
  1337 => (x"66",x"c4",x"4b",x"bf"),
  1338 => (x"12",x"2c",x"73",x"4c"),
  1339 => (x"58",x"a6",x"cc",x"48"),
  1340 => (x"84",x"c1",x"9c",x"70"),
  1341 => (x"69",x"97",x"81",x"c9"),
  1342 => (x"04",x"ac",x"b7",x"49"),
  1343 => (x"4c",x"c0",x"87",x"c2"),
  1344 => (x"4a",x"bf",x"97",x"6e"),
  1345 => (x"72",x"49",x"66",x"c8"),
  1346 => (x"c4",x"b9",x"ff",x"31"),
  1347 => (x"48",x"74",x"99",x"66"),
  1348 => (x"4a",x"70",x"30",x"72"),
  1349 => (x"e4",x"f0",x"c2",x"b1"),
  1350 => (x"f9",x"fd",x"71",x"59"),
  1351 => (x"c2",x"1e",x"c7",x"87"),
  1352 => (x"1e",x"bf",x"c0",x"f1"),
  1353 => (x"1e",x"ec",x"ec",x"c1"),
  1354 => (x"97",x"e4",x"f0",x"c2"),
  1355 => (x"f4",x"c1",x"49",x"bf"),
  1356 => (x"c0",x"49",x"75",x"87"),
  1357 => (x"e8",x"87",x"c9",x"f6"),
  1358 => (x"26",x"4d",x"26",x"8e"),
  1359 => (x"26",x"4b",x"26",x"4c"),
  1360 => (x"1e",x"73",x"1e",x"4f"),
  1361 => (x"fd",x"49",x"4b",x"71"),
  1362 => (x"49",x"73",x"87",x"f9"),
  1363 => (x"26",x"87",x"f4",x"fd"),
  1364 => (x"1e",x"4f",x"26",x"4b"),
  1365 => (x"4b",x"71",x"1e",x"73"),
  1366 => (x"02",x"4a",x"a3",x"c2"),
  1367 => (x"8a",x"c1",x"87",x"d6"),
  1368 => (x"87",x"e2",x"c0",x"05"),
  1369 => (x"bf",x"c0",x"f1",x"c2"),
  1370 => (x"48",x"87",x"db",x"02"),
  1371 => (x"f1",x"c2",x"88",x"c1"),
  1372 => (x"87",x"d2",x"58",x"c4"),
  1373 => (x"bf",x"c4",x"f1",x"c2"),
  1374 => (x"c2",x"87",x"cb",x"02"),
  1375 => (x"48",x"bf",x"c0",x"f1"),
  1376 => (x"f1",x"c2",x"80",x"c1"),
  1377 => (x"1e",x"c7",x"58",x"c4"),
  1378 => (x"bf",x"c0",x"f1",x"c2"),
  1379 => (x"ec",x"ec",x"c1",x"1e"),
  1380 => (x"e4",x"f0",x"c2",x"1e"),
  1381 => (x"cc",x"49",x"bf",x"97"),
  1382 => (x"c0",x"49",x"73",x"87"),
  1383 => (x"f4",x"87",x"e1",x"f4"),
  1384 => (x"26",x"4b",x"26",x"8e"),
  1385 => (x"5b",x"5e",x"0e",x"4f"),
  1386 => (x"ff",x"0e",x"5d",x"5c"),
  1387 => (x"e4",x"c0",x"86",x"cc"),
  1388 => (x"a6",x"cc",x"59",x"a6"),
  1389 => (x"c4",x"78",x"c0",x"48"),
  1390 => (x"c4",x"78",x"c0",x"80"),
  1391 => (x"66",x"c8",x"c1",x"80"),
  1392 => (x"c1",x"80",x"c4",x"78"),
  1393 => (x"c1",x"80",x"c4",x"78"),
  1394 => (x"c4",x"f1",x"c2",x"78"),
  1395 => (x"e0",x"78",x"c1",x"48"),
  1396 => (x"c4",x"e1",x"87",x"ea"),
  1397 => (x"87",x"d9",x"e0",x"87"),
  1398 => (x"fb",x"c0",x"4c",x"70"),
  1399 => (x"f3",x"c1",x"02",x"ac"),
  1400 => (x"66",x"e0",x"c0",x"87"),
  1401 => (x"87",x"e8",x"c1",x"05"),
  1402 => (x"4a",x"66",x"c4",x"c1"),
  1403 => (x"7e",x"6a",x"82",x"c4"),
  1404 => (x"48",x"fc",x"e8",x"c1"),
  1405 => (x"41",x"20",x"49",x"6e"),
  1406 => (x"51",x"10",x"41",x"20"),
  1407 => (x"48",x"66",x"c4",x"c1"),
  1408 => (x"78",x"ef",x"d0",x"c1"),
  1409 => (x"81",x"c7",x"49",x"6a"),
  1410 => (x"c4",x"c1",x"51",x"74"),
  1411 => (x"81",x"c8",x"49",x"66"),
  1412 => (x"a6",x"d8",x"51",x"c1"),
  1413 => (x"c1",x"78",x"c2",x"48"),
  1414 => (x"c9",x"49",x"66",x"c4"),
  1415 => (x"c1",x"51",x"c0",x"81"),
  1416 => (x"ca",x"49",x"66",x"c4"),
  1417 => (x"c1",x"51",x"c0",x"81"),
  1418 => (x"6a",x"1e",x"d8",x"1e"),
  1419 => (x"ff",x"81",x"c8",x"49"),
  1420 => (x"c8",x"87",x"fa",x"df"),
  1421 => (x"66",x"c8",x"c1",x"86"),
  1422 => (x"01",x"a8",x"c0",x"48"),
  1423 => (x"a6",x"d0",x"87",x"c7"),
  1424 => (x"cf",x"78",x"c1",x"48"),
  1425 => (x"66",x"c8",x"c1",x"87"),
  1426 => (x"d8",x"88",x"c1",x"48"),
  1427 => (x"87",x"c4",x"58",x"a6"),
  1428 => (x"87",x"c5",x"df",x"ff"),
  1429 => (x"cd",x"02",x"9c",x"74"),
  1430 => (x"66",x"d0",x"87",x"d9"),
  1431 => (x"66",x"cc",x"c1",x"48"),
  1432 => (x"ce",x"cd",x"03",x"a8"),
  1433 => (x"48",x"a6",x"c8",x"87"),
  1434 => (x"ff",x"7e",x"78",x"c0"),
  1435 => (x"70",x"87",x"c2",x"de"),
  1436 => (x"ac",x"d0",x"c1",x"4c"),
  1437 => (x"87",x"e7",x"c2",x"05"),
  1438 => (x"6e",x"48",x"a6",x"c4"),
  1439 => (x"87",x"d8",x"e0",x"78"),
  1440 => (x"cc",x"48",x"7e",x"70"),
  1441 => (x"c5",x"06",x"a8",x"66"),
  1442 => (x"48",x"a6",x"cc",x"87"),
  1443 => (x"dd",x"ff",x"78",x"6e"),
  1444 => (x"4c",x"70",x"87",x"df"),
  1445 => (x"05",x"ac",x"ec",x"c0"),
  1446 => (x"d0",x"87",x"ee",x"c1"),
  1447 => (x"91",x"cc",x"49",x"66"),
  1448 => (x"81",x"66",x"c4",x"c1"),
  1449 => (x"6a",x"4a",x"a1",x"c4"),
  1450 => (x"4a",x"a1",x"c8",x"4d"),
  1451 => (x"d1",x"c1",x"52",x"6e"),
  1452 => (x"dc",x"ff",x"79",x"f5"),
  1453 => (x"4c",x"70",x"87",x"fb"),
  1454 => (x"87",x"d9",x"02",x"9c"),
  1455 => (x"02",x"ac",x"fb",x"c0"),
  1456 => (x"55",x"74",x"87",x"d3"),
  1457 => (x"87",x"e9",x"dc",x"ff"),
  1458 => (x"02",x"9c",x"4c",x"70"),
  1459 => (x"fb",x"c0",x"87",x"c7"),
  1460 => (x"ed",x"ff",x"05",x"ac"),
  1461 => (x"55",x"e0",x"c0",x"87"),
  1462 => (x"c0",x"55",x"c1",x"c2"),
  1463 => (x"e0",x"c0",x"7d",x"97"),
  1464 => (x"66",x"c4",x"48",x"66"),
  1465 => (x"87",x"db",x"05",x"a8"),
  1466 => (x"d4",x"48",x"66",x"d0"),
  1467 => (x"ca",x"04",x"a8",x"66"),
  1468 => (x"48",x"66",x"d0",x"87"),
  1469 => (x"a6",x"d4",x"80",x"c1"),
  1470 => (x"d4",x"87",x"c8",x"58"),
  1471 => (x"88",x"c1",x"48",x"66"),
  1472 => (x"ff",x"58",x"a6",x"d8"),
  1473 => (x"70",x"87",x"ea",x"db"),
  1474 => (x"ac",x"d0",x"c1",x"4c"),
  1475 => (x"dc",x"87",x"c9",x"05"),
  1476 => (x"80",x"c1",x"48",x"66"),
  1477 => (x"58",x"a6",x"e0",x"c0"),
  1478 => (x"02",x"ac",x"d0",x"c1"),
  1479 => (x"6e",x"87",x"d9",x"fd"),
  1480 => (x"66",x"e0",x"c0",x"48"),
  1481 => (x"ea",x"c9",x"05",x"a8"),
  1482 => (x"a6",x"e4",x"c0",x"87"),
  1483 => (x"74",x"78",x"c0",x"48"),
  1484 => (x"88",x"fb",x"c0",x"48"),
  1485 => (x"70",x"58",x"a6",x"c8"),
  1486 => (x"dc",x"c9",x"02",x"98"),
  1487 => (x"88",x"cb",x"48",x"87"),
  1488 => (x"70",x"58",x"a6",x"c8"),
  1489 => (x"ce",x"c1",x"02",x"98"),
  1490 => (x"88",x"c9",x"48",x"87"),
  1491 => (x"70",x"58",x"a6",x"c8"),
  1492 => (x"fe",x"c3",x"02",x"98"),
  1493 => (x"88",x"c4",x"48",x"87"),
  1494 => (x"70",x"58",x"a6",x"c8"),
  1495 => (x"87",x"cf",x"02",x"98"),
  1496 => (x"c8",x"88",x"c1",x"48"),
  1497 => (x"98",x"70",x"58",x"a6"),
  1498 => (x"87",x"e7",x"c3",x"02"),
  1499 => (x"c8",x"87",x"db",x"c8"),
  1500 => (x"f0",x"c0",x"48",x"a6"),
  1501 => (x"f8",x"d9",x"ff",x"78"),
  1502 => (x"c0",x"4c",x"70",x"87"),
  1503 => (x"c3",x"02",x"ac",x"ec"),
  1504 => (x"5c",x"a6",x"cc",x"87"),
  1505 => (x"02",x"ac",x"ec",x"c0"),
  1506 => (x"d9",x"ff",x"87",x"cd"),
  1507 => (x"4c",x"70",x"87",x"e3"),
  1508 => (x"05",x"ac",x"ec",x"c0"),
  1509 => (x"c0",x"87",x"f3",x"ff"),
  1510 => (x"c0",x"02",x"ac",x"ec"),
  1511 => (x"d9",x"ff",x"87",x"c4"),
  1512 => (x"1e",x"c0",x"87",x"cf"),
  1513 => (x"66",x"d8",x"1e",x"ca"),
  1514 => (x"c1",x"91",x"cc",x"49"),
  1515 => (x"71",x"48",x"66",x"cc"),
  1516 => (x"58",x"a6",x"cc",x"80"),
  1517 => (x"c4",x"48",x"66",x"c8"),
  1518 => (x"58",x"a6",x"d0",x"80"),
  1519 => (x"49",x"bf",x"66",x"cc"),
  1520 => (x"87",x"e9",x"d9",x"ff"),
  1521 => (x"1e",x"de",x"1e",x"c1"),
  1522 => (x"49",x"bf",x"66",x"d4"),
  1523 => (x"87",x"dd",x"d9",x"ff"),
  1524 => (x"49",x"70",x"86",x"d0"),
  1525 => (x"88",x"08",x"c0",x"48"),
  1526 => (x"58",x"a6",x"ec",x"c0"),
  1527 => (x"c0",x"06",x"a8",x"c0"),
  1528 => (x"e8",x"c0",x"87",x"ee"),
  1529 => (x"a8",x"dd",x"48",x"66"),
  1530 => (x"87",x"e4",x"c0",x"03"),
  1531 => (x"49",x"bf",x"66",x"c4"),
  1532 => (x"81",x"66",x"e8",x"c0"),
  1533 => (x"c0",x"51",x"e0",x"c0"),
  1534 => (x"c1",x"49",x"66",x"e8"),
  1535 => (x"bf",x"66",x"c4",x"81"),
  1536 => (x"51",x"c1",x"c2",x"81"),
  1537 => (x"49",x"66",x"e8",x"c0"),
  1538 => (x"66",x"c4",x"81",x"c2"),
  1539 => (x"51",x"c0",x"81",x"bf"),
  1540 => (x"d0",x"c1",x"48",x"6e"),
  1541 => (x"49",x"6e",x"78",x"ef"),
  1542 => (x"66",x"d8",x"81",x"c8"),
  1543 => (x"c9",x"49",x"6e",x"51"),
  1544 => (x"51",x"66",x"dc",x"81"),
  1545 => (x"81",x"ca",x"49",x"6e"),
  1546 => (x"d8",x"51",x"66",x"c8"),
  1547 => (x"80",x"c1",x"48",x"66"),
  1548 => (x"d0",x"58",x"a6",x"dc"),
  1549 => (x"66",x"d4",x"48",x"66"),
  1550 => (x"cb",x"c0",x"04",x"a8"),
  1551 => (x"48",x"66",x"d0",x"87"),
  1552 => (x"a6",x"d4",x"80",x"c1"),
  1553 => (x"87",x"d1",x"c5",x"58"),
  1554 => (x"c1",x"48",x"66",x"d4"),
  1555 => (x"58",x"a6",x"d8",x"88"),
  1556 => (x"ff",x"87",x"c6",x"c5"),
  1557 => (x"c0",x"87",x"c1",x"d9"),
  1558 => (x"ff",x"58",x"a6",x"ec"),
  1559 => (x"c0",x"87",x"f9",x"d8"),
  1560 => (x"c0",x"58",x"a6",x"f0"),
  1561 => (x"c0",x"05",x"a8",x"ec"),
  1562 => (x"48",x"a6",x"87",x"c9"),
  1563 => (x"78",x"66",x"e8",x"c0"),
  1564 => (x"ff",x"87",x"c4",x"c0"),
  1565 => (x"d0",x"87",x"fa",x"d5"),
  1566 => (x"91",x"cc",x"49",x"66"),
  1567 => (x"48",x"66",x"c4",x"c1"),
  1568 => (x"a6",x"c8",x"80",x"71"),
  1569 => (x"4a",x"66",x"c4",x"58"),
  1570 => (x"66",x"c4",x"82",x"c8"),
  1571 => (x"c0",x"81",x"ca",x"49"),
  1572 => (x"c0",x"51",x"66",x"e8"),
  1573 => (x"c1",x"49",x"66",x"ec"),
  1574 => (x"66",x"e8",x"c0",x"81"),
  1575 => (x"71",x"48",x"c1",x"89"),
  1576 => (x"c1",x"49",x"70",x"30"),
  1577 => (x"7a",x"97",x"71",x"89"),
  1578 => (x"bf",x"e0",x"f0",x"c2"),
  1579 => (x"66",x"e8",x"c0",x"49"),
  1580 => (x"4a",x"6a",x"97",x"29"),
  1581 => (x"c0",x"98",x"71",x"48"),
  1582 => (x"c4",x"58",x"a6",x"f4"),
  1583 => (x"80",x"c4",x"48",x"66"),
  1584 => (x"c8",x"58",x"a6",x"cc"),
  1585 => (x"c0",x"4d",x"bf",x"66"),
  1586 => (x"6e",x"48",x"66",x"e0"),
  1587 => (x"c5",x"c0",x"02",x"a8"),
  1588 => (x"c0",x"7e",x"c0",x"87"),
  1589 => (x"7e",x"c1",x"87",x"c2"),
  1590 => (x"e0",x"c0",x"1e",x"6e"),
  1591 => (x"ff",x"49",x"75",x"1e"),
  1592 => (x"c8",x"87",x"ca",x"d5"),
  1593 => (x"c0",x"4c",x"70",x"86"),
  1594 => (x"c1",x"06",x"ac",x"b7"),
  1595 => (x"85",x"74",x"87",x"d4"),
  1596 => (x"49",x"bf",x"66",x"c8"),
  1597 => (x"75",x"81",x"e0",x"c0"),
  1598 => (x"e9",x"c1",x"4b",x"89"),
  1599 => (x"fe",x"71",x"4a",x"c8"),
  1600 => (x"c2",x"87",x"e1",x"e0"),
  1601 => (x"c0",x"7e",x"75",x"85"),
  1602 => (x"c1",x"48",x"66",x"e4"),
  1603 => (x"a6",x"e8",x"c0",x"80"),
  1604 => (x"66",x"f0",x"c0",x"58"),
  1605 => (x"70",x"81",x"c1",x"49"),
  1606 => (x"c5",x"c0",x"02",x"a9"),
  1607 => (x"c0",x"4d",x"c0",x"87"),
  1608 => (x"4d",x"c1",x"87",x"c2"),
  1609 => (x"66",x"cc",x"1e",x"75"),
  1610 => (x"e0",x"c0",x"49",x"bf"),
  1611 => (x"89",x"66",x"c4",x"81"),
  1612 => (x"66",x"c8",x"1e",x"71"),
  1613 => (x"f4",x"d3",x"ff",x"49"),
  1614 => (x"c0",x"86",x"c8",x"87"),
  1615 => (x"ff",x"01",x"a8",x"b7"),
  1616 => (x"e4",x"c0",x"87",x"c5"),
  1617 => (x"d3",x"c0",x"02",x"66"),
  1618 => (x"49",x"66",x"c4",x"87"),
  1619 => (x"e4",x"c0",x"81",x"c9"),
  1620 => (x"66",x"c4",x"51",x"66"),
  1621 => (x"c3",x"d3",x"c1",x"48"),
  1622 => (x"87",x"ce",x"c0",x"78"),
  1623 => (x"c9",x"49",x"66",x"c4"),
  1624 => (x"c4",x"51",x"c2",x"81"),
  1625 => (x"d5",x"c1",x"48",x"66"),
  1626 => (x"66",x"d0",x"78",x"c1"),
  1627 => (x"a8",x"66",x"d4",x"48"),
  1628 => (x"87",x"cb",x"c0",x"04"),
  1629 => (x"c1",x"48",x"66",x"d0"),
  1630 => (x"58",x"a6",x"d4",x"80"),
  1631 => (x"d4",x"87",x"da",x"c0"),
  1632 => (x"88",x"c1",x"48",x"66"),
  1633 => (x"c0",x"58",x"a6",x"d8"),
  1634 => (x"d2",x"ff",x"87",x"cf"),
  1635 => (x"4c",x"70",x"87",x"cb"),
  1636 => (x"ff",x"87",x"c6",x"c0"),
  1637 => (x"70",x"87",x"c2",x"d2"),
  1638 => (x"48",x"66",x"dc",x"4c"),
  1639 => (x"e0",x"c0",x"80",x"c1"),
  1640 => (x"9c",x"74",x"58",x"a6"),
  1641 => (x"87",x"cb",x"c0",x"02"),
  1642 => (x"c1",x"48",x"66",x"d0"),
  1643 => (x"04",x"a8",x"66",x"cc"),
  1644 => (x"d0",x"87",x"f2",x"f2"),
  1645 => (x"a8",x"c7",x"48",x"66"),
  1646 => (x"87",x"e1",x"c0",x"03"),
  1647 => (x"c2",x"4c",x"66",x"d0"),
  1648 => (x"c0",x"48",x"c4",x"f1"),
  1649 => (x"cc",x"49",x"74",x"78"),
  1650 => (x"66",x"c4",x"c1",x"91"),
  1651 => (x"4a",x"a1",x"c4",x"81"),
  1652 => (x"52",x"c0",x"4a",x"6a"),
  1653 => (x"c7",x"84",x"c1",x"79"),
  1654 => (x"e2",x"ff",x"04",x"ac"),
  1655 => (x"66",x"e0",x"c0",x"87"),
  1656 => (x"87",x"e2",x"c0",x"02"),
  1657 => (x"49",x"66",x"c4",x"c1"),
  1658 => (x"c1",x"81",x"d4",x"c1"),
  1659 => (x"c1",x"4a",x"66",x"c4"),
  1660 => (x"52",x"c0",x"82",x"dc"),
  1661 => (x"79",x"f5",x"d1",x"c1"),
  1662 => (x"49",x"66",x"c4",x"c1"),
  1663 => (x"c1",x"81",x"d8",x"c1"),
  1664 => (x"c0",x"79",x"cc",x"e9"),
  1665 => (x"c4",x"c1",x"87",x"d6"),
  1666 => (x"d4",x"c1",x"49",x"66"),
  1667 => (x"66",x"c4",x"c1",x"81"),
  1668 => (x"82",x"d8",x"c1",x"4a"),
  1669 => (x"7a",x"d4",x"e9",x"c1"),
  1670 => (x"79",x"ec",x"d1",x"c1"),
  1671 => (x"49",x"66",x"c4",x"c1"),
  1672 => (x"c1",x"81",x"e0",x"c1"),
  1673 => (x"ff",x"79",x"d3",x"d5"),
  1674 => (x"cc",x"87",x"e5",x"cf"),
  1675 => (x"cc",x"ff",x"48",x"66"),
  1676 => (x"26",x"4d",x"26",x"8e"),
  1677 => (x"26",x"4b",x"26",x"4c"),
  1678 => (x"00",x"00",x"00",x"4f"),
  1679 => (x"64",x"61",x"6f",x"4c"),
  1680 => (x"20",x"2e",x"2a",x"20"),
  1681 => (x"00",x"00",x"00",x"00"),
  1682 => (x"00",x"00",x"20",x"3a"),
  1683 => (x"61",x"42",x"20",x"80"),
  1684 => (x"00",x"00",x"6b",x"63"),
  1685 => (x"78",x"45",x"20",x"80"),
  1686 => (x"1e",x"00",x"74",x"69"),
  1687 => (x"f1",x"c2",x"1e",x"c7"),
  1688 => (x"c1",x"1e",x"bf",x"c0"),
  1689 => (x"c2",x"1e",x"ec",x"ec"),
  1690 => (x"bf",x"97",x"e4",x"f0"),
  1691 => (x"87",x"f5",x"ec",x"49"),
  1692 => (x"49",x"ec",x"ec",x"c1"),
  1693 => (x"87",x"d6",x"e2",x"c0"),
  1694 => (x"4f",x"26",x"8e",x"f4"),
  1695 => (x"c8",x"1e",x"73",x"1e"),
  1696 => (x"ee",x"c1",x"87",x"c3"),
  1697 => (x"ec",x"c1",x"48",x"c4"),
  1698 => (x"e8",x"fe",x"78",x"cc"),
  1699 => (x"e1",x"c0",x"49",x"a0"),
  1700 => (x"49",x"c7",x"87",x"fc"),
  1701 => (x"87",x"e8",x"e0",x"c0"),
  1702 => (x"e2",x"c0",x"49",x"c1"),
  1703 => (x"d4",x"ff",x"87",x"c3"),
  1704 => (x"78",x"ff",x"c3",x"48"),
  1705 => (x"48",x"cc",x"f1",x"c2"),
  1706 => (x"e3",x"fe",x"50",x"c0"),
  1707 => (x"98",x"70",x"87",x"de"),
  1708 => (x"fe",x"87",x"cd",x"02"),
  1709 => (x"70",x"87",x"da",x"ed"),
  1710 => (x"87",x"c4",x"02",x"98"),
  1711 => (x"87",x"c2",x"4a",x"c1"),
  1712 => (x"9a",x"72",x"4a",x"c0"),
  1713 => (x"c1",x"87",x"c8",x"02"),
  1714 => (x"fe",x"49",x"d8",x"ec"),
  1715 => (x"c2",x"87",x"d8",x"d7"),
  1716 => (x"c0",x"48",x"c0",x"f1"),
  1717 => (x"e4",x"f0",x"c2",x"78"),
  1718 => (x"49",x"50",x"c0",x"48"),
  1719 => (x"c0",x"87",x"fc",x"fd"),
  1720 => (x"70",x"87",x"cd",x"f6"),
  1721 => (x"cb",x"02",x"9b",x"4b"),
  1722 => (x"c8",x"ee",x"c1",x"87"),
  1723 => (x"df",x"49",x"c7",x"5b"),
  1724 => (x"87",x"c6",x"87",x"ce"),
  1725 => (x"e0",x"c0",x"49",x"c0"),
  1726 => (x"c2",x"c3",x"87",x"e7"),
  1727 => (x"c8",x"e2",x"c0",x"87"),
  1728 => (x"d4",x"f0",x"c0",x"87"),
  1729 => (x"87",x"f5",x"ff",x"87"),
  1730 => (x"4f",x"26",x"4b",x"26"),
  1731 => (x"74",x"6f",x"6f",x"42"),
  1732 => (x"2e",x"67",x"6e",x"69"),
  1733 => (x"00",x"00",x"2e",x"2e"),
  1734 => (x"4f",x"20",x"44",x"53"),
  1735 => (x"00",x"00",x"00",x"4b"),
  1736 => (x"00",x"00",x"00",x"00"),
  1737 => (x"00",x"00",x"00",x"00"),
  1738 => (x"00",x"00",x"00",x"01"),
  1739 => (x"00",x"00",x"11",x"5a"),
  1740 => (x"00",x"00",x"2c",x"58"),
  1741 => (x"00",x"00",x"00",x"00"),
  1742 => (x"00",x"00",x"11",x"5a"),
  1743 => (x"00",x"00",x"2c",x"76"),
  1744 => (x"00",x"00",x"00",x"00"),
  1745 => (x"00",x"00",x"11",x"5a"),
  1746 => (x"00",x"00",x"2c",x"94"),
  1747 => (x"00",x"00",x"00",x"00"),
  1748 => (x"00",x"00",x"11",x"5a"),
  1749 => (x"00",x"00",x"2c",x"b2"),
  1750 => (x"00",x"00",x"00",x"00"),
  1751 => (x"00",x"00",x"11",x"5a"),
  1752 => (x"00",x"00",x"2c",x"d0"),
  1753 => (x"00",x"00",x"00",x"00"),
  1754 => (x"00",x"00",x"11",x"5a"),
  1755 => (x"00",x"00",x"2c",x"ee"),
  1756 => (x"00",x"00",x"00",x"00"),
  1757 => (x"00",x"00",x"11",x"5a"),
  1758 => (x"00",x"00",x"2d",x"0c"),
  1759 => (x"00",x"00",x"00",x"00"),
  1760 => (x"00",x"00",x"14",x"75"),
  1761 => (x"00",x"00",x"00",x"00"),
  1762 => (x"00",x"00",x"00",x"00"),
  1763 => (x"00",x"00",x"12",x"0f"),
  1764 => (x"00",x"00",x"00",x"00"),
  1765 => (x"00",x"00",x"00",x"00"),
  1766 => (x"db",x"86",x"fc",x"1e"),
  1767 => (x"fc",x"7e",x"70",x"87"),
  1768 => (x"1e",x"4f",x"26",x"8e"),
  1769 => (x"c0",x"48",x"f0",x"fe"),
  1770 => (x"79",x"09",x"cd",x"78"),
  1771 => (x"1e",x"4f",x"26",x"09"),
  1772 => (x"49",x"d8",x"ee",x"c1"),
  1773 => (x"4f",x"26",x"87",x"ed"),
  1774 => (x"bf",x"f0",x"fe",x"1e"),
  1775 => (x"1e",x"4f",x"26",x"48"),
  1776 => (x"c1",x"48",x"f0",x"fe"),
  1777 => (x"1e",x"4f",x"26",x"78"),
  1778 => (x"c0",x"48",x"f0",x"fe"),
  1779 => (x"1e",x"4f",x"26",x"78"),
  1780 => (x"52",x"c0",x"4a",x"71"),
  1781 => (x"0e",x"4f",x"26",x"51"),
  1782 => (x"5d",x"5c",x"5b",x"5e"),
  1783 => (x"71",x"86",x"f4",x"0e"),
  1784 => (x"7e",x"6d",x"97",x"4d"),
  1785 => (x"97",x"4c",x"a5",x"c1"),
  1786 => (x"a6",x"c8",x"48",x"6c"),
  1787 => (x"c4",x"48",x"6e",x"58"),
  1788 => (x"c5",x"05",x"a8",x"66"),
  1789 => (x"c0",x"48",x"ff",x"87"),
  1790 => (x"ca",x"ff",x"87",x"e6"),
  1791 => (x"49",x"a5",x"c2",x"87"),
  1792 => (x"71",x"4b",x"6c",x"97"),
  1793 => (x"6b",x"97",x"4b",x"a3"),
  1794 => (x"7e",x"6c",x"97",x"4b"),
  1795 => (x"80",x"c1",x"48",x"6e"),
  1796 => (x"c7",x"58",x"a6",x"c8"),
  1797 => (x"58",x"a6",x"cc",x"98"),
  1798 => (x"fe",x"7c",x"97",x"70"),
  1799 => (x"48",x"73",x"87",x"e1"),
  1800 => (x"4d",x"26",x"8e",x"f4"),
  1801 => (x"4b",x"26",x"4c",x"26"),
  1802 => (x"5e",x"0e",x"4f",x"26"),
  1803 => (x"f4",x"0e",x"5c",x"5b"),
  1804 => (x"d8",x"4c",x"71",x"86"),
  1805 => (x"ff",x"c3",x"4a",x"66"),
  1806 => (x"4b",x"a4",x"c2",x"9a"),
  1807 => (x"73",x"49",x"6c",x"97"),
  1808 => (x"51",x"72",x"49",x"a1"),
  1809 => (x"6e",x"7e",x"6c",x"97"),
  1810 => (x"c8",x"80",x"c1",x"48"),
  1811 => (x"98",x"c7",x"58",x"a6"),
  1812 => (x"70",x"58",x"a6",x"cc"),
  1813 => (x"26",x"8e",x"f4",x"54"),
  1814 => (x"26",x"4b",x"26",x"4c"),
  1815 => (x"86",x"fc",x"1e",x"4f"),
  1816 => (x"e0",x"87",x"e4",x"fd"),
  1817 => (x"c0",x"49",x"4a",x"bf"),
  1818 => (x"02",x"99",x"c0",x"e0"),
  1819 => (x"1e",x"72",x"87",x"cb"),
  1820 => (x"49",x"ec",x"f4",x"c2"),
  1821 => (x"c4",x"87",x"f3",x"fe"),
  1822 => (x"87",x"fc",x"fc",x"86"),
  1823 => (x"fe",x"fc",x"7e",x"70"),
  1824 => (x"26",x"8e",x"fc",x"87"),
  1825 => (x"f4",x"c2",x"1e",x"4f"),
  1826 => (x"c2",x"fd",x"49",x"ec"),
  1827 => (x"dd",x"f1",x"c1",x"87"),
  1828 => (x"87",x"cf",x"fc",x"49"),
  1829 => (x"26",x"87",x"ed",x"c3"),
  1830 => (x"5b",x"5e",x"0e",x"4f"),
  1831 => (x"fc",x"0e",x"5d",x"5c"),
  1832 => (x"ff",x"7e",x"71",x"86"),
  1833 => (x"f4",x"c2",x"4d",x"d4"),
  1834 => (x"ea",x"fc",x"49",x"ec"),
  1835 => (x"c0",x"4b",x"70",x"87"),
  1836 => (x"c2",x"04",x"ab",x"b7"),
  1837 => (x"f0",x"c3",x"87",x"f8"),
  1838 => (x"87",x"c9",x"05",x"ab"),
  1839 => (x"48",x"fc",x"f5",x"c1"),
  1840 => (x"d9",x"c2",x"78",x"c1"),
  1841 => (x"ab",x"e0",x"c3",x"87"),
  1842 => (x"c1",x"87",x"c9",x"05"),
  1843 => (x"c1",x"48",x"c0",x"f6"),
  1844 => (x"87",x"ca",x"c2",x"78"),
  1845 => (x"bf",x"c0",x"f6",x"c1"),
  1846 => (x"c2",x"87",x"c6",x"02"),
  1847 => (x"c2",x"4c",x"a3",x"c0"),
  1848 => (x"c1",x"4c",x"73",x"87"),
  1849 => (x"02",x"bf",x"fc",x"f5"),
  1850 => (x"74",x"87",x"e0",x"c0"),
  1851 => (x"29",x"b7",x"c4",x"49"),
  1852 => (x"d8",x"f7",x"c1",x"91"),
  1853 => (x"cf",x"4a",x"74",x"81"),
  1854 => (x"c1",x"92",x"c2",x"9a"),
  1855 => (x"70",x"30",x"72",x"48"),
  1856 => (x"72",x"ba",x"ff",x"4a"),
  1857 => (x"70",x"98",x"69",x"48"),
  1858 => (x"74",x"87",x"db",x"79"),
  1859 => (x"29",x"b7",x"c4",x"49"),
  1860 => (x"d8",x"f7",x"c1",x"91"),
  1861 => (x"cf",x"4a",x"74",x"81"),
  1862 => (x"c3",x"92",x"c2",x"9a"),
  1863 => (x"70",x"30",x"72",x"48"),
  1864 => (x"b0",x"69",x"48",x"4a"),
  1865 => (x"05",x"6e",x"79",x"70"),
  1866 => (x"ff",x"87",x"e7",x"c0"),
  1867 => (x"e1",x"c8",x"48",x"d0"),
  1868 => (x"c1",x"7d",x"c5",x"78"),
  1869 => (x"02",x"bf",x"c0",x"f6"),
  1870 => (x"e0",x"c3",x"87",x"c3"),
  1871 => (x"fc",x"f5",x"c1",x"7d"),
  1872 => (x"87",x"c3",x"02",x"bf"),
  1873 => (x"73",x"7d",x"f0",x"c3"),
  1874 => (x"48",x"d0",x"ff",x"7d"),
  1875 => (x"c0",x"78",x"e1",x"c8"),
  1876 => (x"f6",x"c1",x"78",x"e0"),
  1877 => (x"78",x"c0",x"48",x"c0"),
  1878 => (x"48",x"fc",x"f5",x"c1"),
  1879 => (x"f4",x"c2",x"78",x"c0"),
  1880 => (x"f2",x"f9",x"49",x"ec"),
  1881 => (x"c0",x"4b",x"70",x"87"),
  1882 => (x"fd",x"03",x"ab",x"b7"),
  1883 => (x"48",x"c0",x"87",x"c8"),
  1884 => (x"4d",x"26",x"8e",x"fc"),
  1885 => (x"4b",x"26",x"4c",x"26"),
  1886 => (x"00",x"00",x"4f",x"26"),
  1887 => (x"00",x"00",x"00",x"00"),
  1888 => (x"00",x"00",x"00",x"00"),
  1889 => (x"72",x"4a",x"c0",x"1e"),
  1890 => (x"c1",x"91",x"c4",x"49"),
  1891 => (x"c0",x"81",x"d8",x"f7"),
  1892 => (x"d0",x"82",x"c1",x"79"),
  1893 => (x"ee",x"04",x"aa",x"b7"),
  1894 => (x"0e",x"4f",x"26",x"87"),
  1895 => (x"5d",x"5c",x"5b",x"5e"),
  1896 => (x"f8",x"4d",x"71",x"0e"),
  1897 => (x"4a",x"75",x"87",x"e1"),
  1898 => (x"92",x"2a",x"b7",x"c4"),
  1899 => (x"82",x"d8",x"f7",x"c1"),
  1900 => (x"9c",x"cf",x"4c",x"75"),
  1901 => (x"49",x"6a",x"94",x"c2"),
  1902 => (x"c3",x"2b",x"74",x"4b"),
  1903 => (x"74",x"48",x"c2",x"9b"),
  1904 => (x"ff",x"4c",x"70",x"30"),
  1905 => (x"71",x"48",x"74",x"bc"),
  1906 => (x"f7",x"7a",x"70",x"98"),
  1907 => (x"48",x"73",x"87",x"f1"),
  1908 => (x"4c",x"26",x"4d",x"26"),
  1909 => (x"4f",x"26",x"4b",x"26"),
  1910 => (x"00",x"00",x"00",x"00"),
  1911 => (x"00",x"00",x"00",x"00"),
  1912 => (x"00",x"00",x"00",x"00"),
  1913 => (x"00",x"00",x"00",x"00"),
  1914 => (x"00",x"00",x"00",x"00"),
  1915 => (x"00",x"00",x"00",x"00"),
  1916 => (x"00",x"00",x"00",x"00"),
  1917 => (x"00",x"00",x"00",x"00"),
  1918 => (x"00",x"00",x"00",x"00"),
  1919 => (x"00",x"00",x"00",x"00"),
  1920 => (x"00",x"00",x"00",x"00"),
  1921 => (x"00",x"00",x"00",x"00"),
  1922 => (x"00",x"00",x"00",x"00"),
  1923 => (x"00",x"00",x"00",x"00"),
  1924 => (x"00",x"00",x"00",x"00"),
  1925 => (x"00",x"00",x"00",x"00"),
  1926 => (x"48",x"d0",x"ff",x"1e"),
  1927 => (x"71",x"78",x"e1",x"c8"),
  1928 => (x"08",x"d4",x"ff",x"48"),
  1929 => (x"1e",x"4f",x"26",x"78"),
  1930 => (x"c8",x"48",x"d0",x"ff"),
  1931 => (x"48",x"71",x"78",x"e1"),
  1932 => (x"78",x"08",x"d4",x"ff"),
  1933 => (x"ff",x"48",x"66",x"c4"),
  1934 => (x"26",x"78",x"08",x"d4"),
  1935 => (x"4a",x"71",x"1e",x"4f"),
  1936 => (x"1e",x"49",x"66",x"c4"),
  1937 => (x"de",x"ff",x"49",x"72"),
  1938 => (x"48",x"d0",x"ff",x"87"),
  1939 => (x"fc",x"78",x"e0",x"c0"),
  1940 => (x"1e",x"4f",x"26",x"8e"),
  1941 => (x"4b",x"71",x"1e",x"73"),
  1942 => (x"1e",x"49",x"66",x"c8"),
  1943 => (x"e0",x"c1",x"4a",x"73"),
  1944 => (x"d8",x"ff",x"49",x"a2"),
  1945 => (x"26",x"8e",x"fc",x"87"),
  1946 => (x"1e",x"4f",x"26",x"4b"),
  1947 => (x"c8",x"48",x"d0",x"ff"),
  1948 => (x"48",x"71",x"78",x"c9"),
  1949 => (x"78",x"08",x"d4",x"ff"),
  1950 => (x"71",x"1e",x"4f",x"26"),
  1951 => (x"87",x"eb",x"49",x"4a"),
  1952 => (x"c8",x"48",x"d0",x"ff"),
  1953 => (x"1e",x"4f",x"26",x"78"),
  1954 => (x"4b",x"71",x"1e",x"73"),
  1955 => (x"bf",x"c4",x"f5",x"c2"),
  1956 => (x"c2",x"87",x"c3",x"02"),
  1957 => (x"d0",x"ff",x"87",x"eb"),
  1958 => (x"78",x"c9",x"c8",x"48"),
  1959 => (x"e0",x"c0",x"48",x"73"),
  1960 => (x"08",x"d4",x"ff",x"b0"),
  1961 => (x"f8",x"f4",x"c2",x"78"),
  1962 => (x"c8",x"78",x"c0",x"48"),
  1963 => (x"87",x"c5",x"02",x"66"),
  1964 => (x"c2",x"49",x"ff",x"c3"),
  1965 => (x"c2",x"49",x"c0",x"87"),
  1966 => (x"cc",x"59",x"c0",x"f5"),
  1967 => (x"87",x"c6",x"02",x"66"),
  1968 => (x"4a",x"d5",x"d5",x"c5"),
  1969 => (x"ff",x"cf",x"87",x"c4"),
  1970 => (x"f5",x"c2",x"4a",x"ff"),
  1971 => (x"f5",x"c2",x"5a",x"c4"),
  1972 => (x"78",x"c1",x"48",x"c4"),
  1973 => (x"4f",x"26",x"4b",x"26"),
  1974 => (x"5c",x"5b",x"5e",x"0e"),
  1975 => (x"4d",x"71",x"0e",x"5d"),
  1976 => (x"bf",x"c0",x"f5",x"c2"),
  1977 => (x"02",x"9d",x"75",x"4b"),
  1978 => (x"c8",x"49",x"87",x"cb"),
  1979 => (x"c0",x"fa",x"c1",x"91"),
  1980 => (x"c4",x"82",x"71",x"4a"),
  1981 => (x"c0",x"fe",x"c1",x"87"),
  1982 => (x"12",x"4c",x"c0",x"4a"),
  1983 => (x"c2",x"99",x"73",x"49"),
  1984 => (x"48",x"bf",x"fc",x"f4"),
  1985 => (x"d4",x"ff",x"b8",x"71"),
  1986 => (x"b7",x"c1",x"78",x"08"),
  1987 => (x"b7",x"c8",x"84",x"2b"),
  1988 => (x"87",x"e7",x"04",x"ac"),
  1989 => (x"bf",x"f8",x"f4",x"c2"),
  1990 => (x"c2",x"80",x"c8",x"48"),
  1991 => (x"26",x"58",x"fc",x"f4"),
  1992 => (x"26",x"4c",x"26",x"4d"),
  1993 => (x"1e",x"4f",x"26",x"4b"),
  1994 => (x"4b",x"71",x"1e",x"73"),
  1995 => (x"02",x"9a",x"4a",x"13"),
  1996 => (x"49",x"72",x"87",x"cb"),
  1997 => (x"13",x"87",x"e1",x"fe"),
  1998 => (x"f5",x"05",x"9a",x"4a"),
  1999 => (x"26",x"4b",x"26",x"87"),
  2000 => (x"f4",x"c2",x"1e",x"4f"),
  2001 => (x"c2",x"49",x"bf",x"f8"),
  2002 => (x"c1",x"48",x"f8",x"f4"),
  2003 => (x"c0",x"c4",x"78",x"a1"),
  2004 => (x"db",x"03",x"a9",x"b7"),
  2005 => (x"48",x"d4",x"ff",x"87"),
  2006 => (x"bf",x"fc",x"f4",x"c2"),
  2007 => (x"f8",x"f4",x"c2",x"78"),
  2008 => (x"f4",x"c2",x"49",x"bf"),
  2009 => (x"a1",x"c1",x"48",x"f8"),
  2010 => (x"b7",x"c0",x"c4",x"78"),
  2011 => (x"87",x"e5",x"04",x"a9"),
  2012 => (x"c8",x"48",x"d0",x"ff"),
  2013 => (x"c4",x"f5",x"c2",x"78"),
  2014 => (x"26",x"78",x"c0",x"48"),
  2015 => (x"00",x"00",x"00",x"4f"),
  2016 => (x"00",x"00",x"00",x"00"),
  2017 => (x"00",x"00",x"00",x"00"),
  2018 => (x"5f",x"00",x"00",x"00"),
  2019 => (x"00",x"00",x"00",x"5f"),
  2020 => (x"00",x"03",x"03",x"00"),
  2021 => (x"00",x"00",x"03",x"03"),
  2022 => (x"14",x"7f",x"7f",x"14"),
  2023 => (x"00",x"14",x"7f",x"7f"),
  2024 => (x"6b",x"2e",x"24",x"00"),
  2025 => (x"00",x"12",x"3a",x"6b"),
  2026 => (x"18",x"36",x"6a",x"4c"),
  2027 => (x"00",x"32",x"56",x"6c"),
  2028 => (x"59",x"4f",x"7e",x"30"),
  2029 => (x"40",x"68",x"3a",x"77"),
  2030 => (x"07",x"04",x"00",x"00"),
  2031 => (x"00",x"00",x"00",x"03"),
  2032 => (x"3e",x"1c",x"00",x"00"),
  2033 => (x"00",x"00",x"41",x"63"),
  2034 => (x"63",x"41",x"00",x"00"),
  2035 => (x"00",x"00",x"1c",x"3e"),
  2036 => (x"1c",x"3e",x"2a",x"08"),
  2037 => (x"08",x"2a",x"3e",x"1c"),
  2038 => (x"3e",x"08",x"08",x"00"),
  2039 => (x"00",x"08",x"08",x"3e"),
  2040 => (x"e0",x"80",x"00",x"00"),
  2041 => (x"00",x"00",x"00",x"60"),
  2042 => (x"08",x"08",x"08",x"00"),
  2043 => (x"00",x"08",x"08",x"08"),
  2044 => (x"60",x"00",x"00",x"00"),
  2045 => (x"00",x"00",x"00",x"60"),
  2046 => (x"18",x"30",x"60",x"40"),
  2047 => (x"01",x"03",x"06",x"0c"),
  2048 => (x"59",x"7f",x"3e",x"00"),
  2049 => (x"00",x"3e",x"7f",x"4d"),
  2050 => (x"7f",x"06",x"04",x"00"),
  2051 => (x"00",x"00",x"00",x"7f"),
  2052 => (x"71",x"63",x"42",x"00"),
  2053 => (x"00",x"46",x"4f",x"59"),
  2054 => (x"49",x"63",x"22",x"00"),
  2055 => (x"00",x"36",x"7f",x"49"),
  2056 => (x"13",x"16",x"1c",x"18"),
  2057 => (x"00",x"10",x"7f",x"7f"),
  2058 => (x"45",x"67",x"27",x"00"),
  2059 => (x"00",x"39",x"7d",x"45"),
  2060 => (x"4b",x"7e",x"3c",x"00"),
  2061 => (x"00",x"30",x"79",x"49"),
  2062 => (x"71",x"01",x"01",x"00"),
  2063 => (x"00",x"07",x"0f",x"79"),
  2064 => (x"49",x"7f",x"36",x"00"),
  2065 => (x"00",x"36",x"7f",x"49"),
  2066 => (x"49",x"4f",x"06",x"00"),
  2067 => (x"00",x"1e",x"3f",x"69"),
  2068 => (x"66",x"00",x"00",x"00"),
  2069 => (x"00",x"00",x"00",x"66"),
  2070 => (x"e6",x"80",x"00",x"00"),
  2071 => (x"00",x"00",x"00",x"66"),
  2072 => (x"14",x"08",x"08",x"00"),
  2073 => (x"00",x"22",x"22",x"14"),
  2074 => (x"14",x"14",x"14",x"00"),
  2075 => (x"00",x"14",x"14",x"14"),
  2076 => (x"14",x"22",x"22",x"00"),
  2077 => (x"00",x"08",x"08",x"14"),
  2078 => (x"51",x"03",x"02",x"00"),
  2079 => (x"00",x"06",x"0f",x"59"),
  2080 => (x"5d",x"41",x"7f",x"3e"),
  2081 => (x"00",x"1e",x"1f",x"55"),
  2082 => (x"09",x"7f",x"7e",x"00"),
  2083 => (x"00",x"7e",x"7f",x"09"),
  2084 => (x"49",x"7f",x"7f",x"00"),
  2085 => (x"00",x"36",x"7f",x"49"),
  2086 => (x"63",x"3e",x"1c",x"00"),
  2087 => (x"00",x"41",x"41",x"41"),
  2088 => (x"41",x"7f",x"7f",x"00"),
  2089 => (x"00",x"1c",x"3e",x"63"),
  2090 => (x"49",x"7f",x"7f",x"00"),
  2091 => (x"00",x"41",x"41",x"49"),
  2092 => (x"09",x"7f",x"7f",x"00"),
  2093 => (x"00",x"01",x"01",x"09"),
  2094 => (x"41",x"7f",x"3e",x"00"),
  2095 => (x"00",x"7a",x"7b",x"49"),
  2096 => (x"08",x"7f",x"7f",x"00"),
  2097 => (x"00",x"7f",x"7f",x"08"),
  2098 => (x"7f",x"41",x"00",x"00"),
  2099 => (x"00",x"00",x"41",x"7f"),
  2100 => (x"40",x"60",x"20",x"00"),
  2101 => (x"00",x"3f",x"7f",x"40"),
  2102 => (x"1c",x"08",x"7f",x"7f"),
  2103 => (x"00",x"41",x"63",x"36"),
  2104 => (x"40",x"7f",x"7f",x"00"),
  2105 => (x"00",x"40",x"40",x"40"),
  2106 => (x"0c",x"06",x"7f",x"7f"),
  2107 => (x"00",x"7f",x"7f",x"06"),
  2108 => (x"0c",x"06",x"7f",x"7f"),
  2109 => (x"00",x"7f",x"7f",x"18"),
  2110 => (x"41",x"7f",x"3e",x"00"),
  2111 => (x"00",x"3e",x"7f",x"41"),
  2112 => (x"09",x"7f",x"7f",x"00"),
  2113 => (x"00",x"06",x"0f",x"09"),
  2114 => (x"61",x"41",x"7f",x"3e"),
  2115 => (x"00",x"40",x"7e",x"7f"),
  2116 => (x"09",x"7f",x"7f",x"00"),
  2117 => (x"00",x"66",x"7f",x"19"),
  2118 => (x"4d",x"6f",x"26",x"00"),
  2119 => (x"00",x"32",x"7b",x"59"),
  2120 => (x"7f",x"01",x"01",x"00"),
  2121 => (x"00",x"01",x"01",x"7f"),
  2122 => (x"40",x"7f",x"3f",x"00"),
  2123 => (x"00",x"3f",x"7f",x"40"),
  2124 => (x"70",x"3f",x"0f",x"00"),
  2125 => (x"00",x"0f",x"3f",x"70"),
  2126 => (x"18",x"30",x"7f",x"7f"),
  2127 => (x"00",x"7f",x"7f",x"30"),
  2128 => (x"1c",x"36",x"63",x"41"),
  2129 => (x"41",x"63",x"36",x"1c"),
  2130 => (x"7c",x"06",x"03",x"01"),
  2131 => (x"01",x"03",x"06",x"7c"),
  2132 => (x"4d",x"59",x"71",x"61"),
  2133 => (x"00",x"41",x"43",x"47"),
  2134 => (x"7f",x"7f",x"00",x"00"),
  2135 => (x"00",x"00",x"41",x"41"),
  2136 => (x"0c",x"06",x"03",x"01"),
  2137 => (x"40",x"60",x"30",x"18"),
  2138 => (x"41",x"41",x"00",x"00"),
  2139 => (x"00",x"00",x"7f",x"7f"),
  2140 => (x"03",x"06",x"0c",x"08"),
  2141 => (x"00",x"08",x"0c",x"06"),
  2142 => (x"80",x"80",x"80",x"80"),
  2143 => (x"00",x"80",x"80",x"80"),
  2144 => (x"03",x"00",x"00",x"00"),
  2145 => (x"00",x"00",x"04",x"07"),
  2146 => (x"54",x"74",x"20",x"00"),
  2147 => (x"00",x"78",x"7c",x"54"),
  2148 => (x"44",x"7f",x"7f",x"00"),
  2149 => (x"00",x"38",x"7c",x"44"),
  2150 => (x"44",x"7c",x"38",x"00"),
  2151 => (x"00",x"00",x"44",x"44"),
  2152 => (x"44",x"7c",x"38",x"00"),
  2153 => (x"00",x"7f",x"7f",x"44"),
  2154 => (x"54",x"7c",x"38",x"00"),
  2155 => (x"00",x"18",x"5c",x"54"),
  2156 => (x"7f",x"7e",x"04",x"00"),
  2157 => (x"00",x"00",x"05",x"05"),
  2158 => (x"a4",x"bc",x"18",x"00"),
  2159 => (x"00",x"7c",x"fc",x"a4"),
  2160 => (x"04",x"7f",x"7f",x"00"),
  2161 => (x"00",x"78",x"7c",x"04"),
  2162 => (x"3d",x"00",x"00",x"00"),
  2163 => (x"00",x"00",x"40",x"7d"),
  2164 => (x"80",x"80",x"80",x"00"),
  2165 => (x"00",x"00",x"7d",x"fd"),
  2166 => (x"10",x"7f",x"7f",x"00"),
  2167 => (x"00",x"44",x"6c",x"38"),
  2168 => (x"3f",x"00",x"00",x"00"),
  2169 => (x"00",x"00",x"40",x"7f"),
  2170 => (x"18",x"0c",x"7c",x"7c"),
  2171 => (x"00",x"78",x"7c",x"0c"),
  2172 => (x"04",x"7c",x"7c",x"00"),
  2173 => (x"00",x"78",x"7c",x"04"),
  2174 => (x"44",x"7c",x"38",x"00"),
  2175 => (x"00",x"38",x"7c",x"44"),
  2176 => (x"24",x"fc",x"fc",x"00"),
  2177 => (x"00",x"18",x"3c",x"24"),
  2178 => (x"24",x"3c",x"18",x"00"),
  2179 => (x"00",x"fc",x"fc",x"24"),
  2180 => (x"04",x"7c",x"7c",x"00"),
  2181 => (x"00",x"08",x"0c",x"04"),
  2182 => (x"54",x"5c",x"48",x"00"),
  2183 => (x"00",x"20",x"74",x"54"),
  2184 => (x"7f",x"3f",x"04",x"00"),
  2185 => (x"00",x"00",x"44",x"44"),
  2186 => (x"40",x"7c",x"3c",x"00"),
  2187 => (x"00",x"7c",x"7c",x"40"),
  2188 => (x"60",x"3c",x"1c",x"00"),
  2189 => (x"00",x"1c",x"3c",x"60"),
  2190 => (x"30",x"60",x"7c",x"3c"),
  2191 => (x"00",x"3c",x"7c",x"60"),
  2192 => (x"10",x"38",x"6c",x"44"),
  2193 => (x"00",x"44",x"6c",x"38"),
  2194 => (x"e0",x"bc",x"1c",x"00"),
  2195 => (x"00",x"1c",x"3c",x"60"),
  2196 => (x"74",x"64",x"44",x"00"),
  2197 => (x"00",x"44",x"4c",x"5c"),
  2198 => (x"3e",x"08",x"08",x"00"),
  2199 => (x"00",x"41",x"41",x"77"),
  2200 => (x"7f",x"00",x"00",x"00"),
  2201 => (x"00",x"00",x"00",x"7f"),
  2202 => (x"77",x"41",x"41",x"00"),
  2203 => (x"00",x"08",x"08",x"3e"),
  2204 => (x"03",x"01",x"01",x"02"),
  2205 => (x"00",x"01",x"02",x"02"),
  2206 => (x"7f",x"7f",x"7f",x"7f"),
  2207 => (x"00",x"7f",x"7f",x"7f"),
  2208 => (x"1c",x"1c",x"08",x"08"),
  2209 => (x"7f",x"7f",x"3e",x"3e"),
  2210 => (x"3e",x"3e",x"7f",x"7f"),
  2211 => (x"08",x"08",x"1c",x"1c"),
  2212 => (x"7c",x"18",x"10",x"00"),
  2213 => (x"00",x"10",x"18",x"7c"),
  2214 => (x"7c",x"30",x"10",x"00"),
  2215 => (x"00",x"10",x"30",x"7c"),
  2216 => (x"60",x"60",x"30",x"10"),
  2217 => (x"00",x"06",x"1e",x"78"),
  2218 => (x"18",x"3c",x"66",x"42"),
  2219 => (x"00",x"42",x"66",x"3c"),
  2220 => (x"c2",x"6a",x"38",x"78"),
  2221 => (x"00",x"38",x"6c",x"c6"),
  2222 => (x"60",x"00",x"00",x"60"),
  2223 => (x"00",x"60",x"00",x"00"),
  2224 => (x"5c",x"5b",x"5e",x"0e"),
  2225 => (x"86",x"fc",x"0e",x"5d"),
  2226 => (x"f5",x"c2",x"7e",x"71"),
  2227 => (x"c0",x"4c",x"bf",x"cc"),
  2228 => (x"c4",x"1e",x"c0",x"4b"),
  2229 => (x"c4",x"02",x"ab",x"66"),
  2230 => (x"c2",x"4d",x"c0",x"87"),
  2231 => (x"75",x"4d",x"c1",x"87"),
  2232 => (x"ee",x"49",x"73",x"1e"),
  2233 => (x"86",x"c8",x"87",x"e1"),
  2234 => (x"ef",x"49",x"e0",x"c0"),
  2235 => (x"a4",x"c4",x"87",x"ea"),
  2236 => (x"f0",x"49",x"6a",x"4a"),
  2237 => (x"c8",x"f1",x"87",x"f1"),
  2238 => (x"c1",x"84",x"cc",x"87"),
  2239 => (x"ab",x"b7",x"c8",x"83"),
  2240 => (x"87",x"cd",x"ff",x"04"),
  2241 => (x"4d",x"26",x"8e",x"fc"),
  2242 => (x"4b",x"26",x"4c",x"26"),
  2243 => (x"71",x"1e",x"4f",x"26"),
  2244 => (x"d0",x"f5",x"c2",x"4a"),
  2245 => (x"d0",x"f5",x"c2",x"5a"),
  2246 => (x"49",x"78",x"c7",x"48"),
  2247 => (x"26",x"87",x"e1",x"fe"),
  2248 => (x"1e",x"73",x"1e",x"4f"),
  2249 => (x"b7",x"c0",x"4a",x"71"),
  2250 => (x"87",x"d3",x"03",x"aa"),
  2251 => (x"bf",x"fc",x"d9",x"c2"),
  2252 => (x"c1",x"87",x"c4",x"05"),
  2253 => (x"c0",x"87",x"c2",x"4b"),
  2254 => (x"c0",x"da",x"c2",x"4b"),
  2255 => (x"c2",x"87",x"c4",x"5b"),
  2256 => (x"fc",x"5a",x"c0",x"da"),
  2257 => (x"fc",x"d9",x"c2",x"48"),
  2258 => (x"c1",x"4a",x"78",x"bf"),
  2259 => (x"a2",x"c0",x"c1",x"9a"),
  2260 => (x"87",x"e6",x"ec",x"49"),
  2261 => (x"4f",x"26",x"4b",x"26"),
  2262 => (x"c4",x"4a",x"71",x"1e"),
  2263 => (x"49",x"72",x"1e",x"66"),
  2264 => (x"fc",x"87",x"f0",x"eb"),
  2265 => (x"1e",x"4f",x"26",x"8e"),
  2266 => (x"c3",x"48",x"d4",x"ff"),
  2267 => (x"d0",x"ff",x"78",x"ff"),
  2268 => (x"78",x"e1",x"c0",x"48"),
  2269 => (x"c1",x"48",x"d4",x"ff"),
  2270 => (x"c4",x"48",x"71",x"78"),
  2271 => (x"08",x"d4",x"ff",x"30"),
  2272 => (x"48",x"d0",x"ff",x"78"),
  2273 => (x"26",x"78",x"e0",x"c0"),
  2274 => (x"5b",x"5e",x"0e",x"4f"),
  2275 => (x"ec",x"0e",x"5d",x"5c"),
  2276 => (x"48",x"a6",x"c8",x"86"),
  2277 => (x"c4",x"7e",x"78",x"c0"),
  2278 => (x"78",x"bf",x"ec",x"80"),
  2279 => (x"f5",x"c2",x"80",x"f8"),
  2280 => (x"e8",x"78",x"bf",x"cc"),
  2281 => (x"d9",x"c2",x"4c",x"bf"),
  2282 => (x"e3",x"49",x"bf",x"fc"),
  2283 => (x"ee",x"cb",x"87",x"eb"),
  2284 => (x"87",x"cc",x"cb",x"49"),
  2285 => (x"c7",x"58",x"a6",x"d4"),
  2286 => (x"87",x"df",x"e7",x"49"),
  2287 => (x"c9",x"05",x"98",x"70"),
  2288 => (x"49",x"66",x"cc",x"87"),
  2289 => (x"c1",x"02",x"99",x"c1"),
  2290 => (x"66",x"d0",x"87",x"c4"),
  2291 => (x"ec",x"7e",x"c1",x"4d"),
  2292 => (x"d9",x"c2",x"4b",x"bf"),
  2293 => (x"e2",x"49",x"bf",x"fc"),
  2294 => (x"49",x"75",x"87",x"ff"),
  2295 => (x"70",x"87",x"ed",x"ca"),
  2296 => (x"87",x"d7",x"02",x"98"),
  2297 => (x"bf",x"e4",x"d9",x"c2"),
  2298 => (x"c2",x"b9",x"c1",x"49"),
  2299 => (x"71",x"59",x"e8",x"d9"),
  2300 => (x"cb",x"87",x"f4",x"fd"),
  2301 => (x"c7",x"ca",x"49",x"ee"),
  2302 => (x"c7",x"4d",x"70",x"87"),
  2303 => (x"87",x"db",x"e6",x"49"),
  2304 => (x"ff",x"05",x"98",x"70"),
  2305 => (x"49",x"73",x"87",x"c7"),
  2306 => (x"fe",x"05",x"99",x"c1"),
  2307 => (x"02",x"6e",x"87",x"ff"),
  2308 => (x"c2",x"87",x"e3",x"c0"),
  2309 => (x"4a",x"bf",x"fc",x"d9"),
  2310 => (x"da",x"c2",x"ba",x"c1"),
  2311 => (x"0a",x"fc",x"5a",x"c0"),
  2312 => (x"9a",x"c1",x"0a",x"7a"),
  2313 => (x"49",x"a2",x"c0",x"c1"),
  2314 => (x"c1",x"87",x"cf",x"e9"),
  2315 => (x"ea",x"e5",x"49",x"da"),
  2316 => (x"48",x"a6",x"c8",x"87"),
  2317 => (x"d9",x"c2",x"78",x"c1"),
  2318 => (x"c1",x"05",x"bf",x"fc"),
  2319 => (x"c0",x"c8",x"87",x"c5"),
  2320 => (x"d9",x"c2",x"4d",x"c0"),
  2321 => (x"49",x"13",x"4b",x"e8"),
  2322 => (x"87",x"cf",x"e5",x"49"),
  2323 => (x"c2",x"02",x"98",x"70"),
  2324 => (x"c1",x"b4",x"75",x"87"),
  2325 => (x"ff",x"05",x"2d",x"b7"),
  2326 => (x"49",x"74",x"87",x"ec"),
  2327 => (x"71",x"99",x"ff",x"c3"),
  2328 => (x"fb",x"49",x"c0",x"1e"),
  2329 => (x"49",x"74",x"87",x"f2"),
  2330 => (x"71",x"29",x"b7",x"c8"),
  2331 => (x"fb",x"49",x"c1",x"1e"),
  2332 => (x"86",x"c8",x"87",x"e6"),
  2333 => (x"e4",x"49",x"fd",x"c3"),
  2334 => (x"fa",x"c3",x"87",x"e1"),
  2335 => (x"87",x"db",x"e4",x"49"),
  2336 => (x"74",x"87",x"d4",x"c7"),
  2337 => (x"99",x"ff",x"c3",x"49"),
  2338 => (x"71",x"2c",x"b7",x"c8"),
  2339 => (x"02",x"9c",x"74",x"b4"),
  2340 => (x"d9",x"c2",x"87",x"df"),
  2341 => (x"c7",x"49",x"bf",x"f8"),
  2342 => (x"98",x"70",x"87",x"f2"),
  2343 => (x"87",x"c4",x"c0",x"05"),
  2344 => (x"87",x"d3",x"4c",x"c0"),
  2345 => (x"c7",x"49",x"e0",x"c2"),
  2346 => (x"d9",x"c2",x"87",x"d6"),
  2347 => (x"c6",x"c0",x"58",x"fc"),
  2348 => (x"f8",x"d9",x"c2",x"87"),
  2349 => (x"74",x"78",x"c0",x"48"),
  2350 => (x"05",x"99",x"c8",x"49"),
  2351 => (x"c3",x"87",x"ce",x"c0"),
  2352 => (x"d6",x"e3",x"49",x"f5"),
  2353 => (x"c2",x"49",x"70",x"87"),
  2354 => (x"e7",x"c0",x"02",x"99"),
  2355 => (x"d0",x"f5",x"c2",x"87"),
  2356 => (x"ca",x"c0",x"02",x"bf"),
  2357 => (x"88",x"c1",x"48",x"87"),
  2358 => (x"58",x"d4",x"f5",x"c2"),
  2359 => (x"c4",x"87",x"d0",x"c0"),
  2360 => (x"e0",x"c1",x"4a",x"66"),
  2361 => (x"c0",x"02",x"6a",x"82"),
  2362 => (x"ff",x"4b",x"87",x"c5"),
  2363 => (x"c8",x"0f",x"73",x"49"),
  2364 => (x"78",x"c1",x"48",x"a6"),
  2365 => (x"99",x"c4",x"49",x"74"),
  2366 => (x"87",x"ce",x"c0",x"05"),
  2367 => (x"e2",x"49",x"f2",x"c3"),
  2368 => (x"49",x"70",x"87",x"d9"),
  2369 => (x"c0",x"02",x"99",x"c2"),
  2370 => (x"f5",x"c2",x"87",x"f0"),
  2371 => (x"48",x"7e",x"bf",x"d0"),
  2372 => (x"03",x"a8",x"b7",x"c7"),
  2373 => (x"6e",x"87",x"cb",x"c0"),
  2374 => (x"c2",x"80",x"c1",x"48"),
  2375 => (x"c0",x"58",x"d4",x"f5"),
  2376 => (x"66",x"c4",x"87",x"d3"),
  2377 => (x"80",x"e0",x"c1",x"48"),
  2378 => (x"bf",x"6e",x"7e",x"70"),
  2379 => (x"87",x"c5",x"c0",x"02"),
  2380 => (x"73",x"49",x"fe",x"4b"),
  2381 => (x"48",x"a6",x"c8",x"0f"),
  2382 => (x"fd",x"c3",x"78",x"c1"),
  2383 => (x"87",x"db",x"e1",x"49"),
  2384 => (x"99",x"c2",x"49",x"70"),
  2385 => (x"87",x"e9",x"c0",x"02"),
  2386 => (x"bf",x"d0",x"f5",x"c2"),
  2387 => (x"87",x"c9",x"c0",x"02"),
  2388 => (x"48",x"d0",x"f5",x"c2"),
  2389 => (x"d3",x"c0",x"78",x"c0"),
  2390 => (x"48",x"66",x"c4",x"87"),
  2391 => (x"70",x"80",x"e0",x"c1"),
  2392 => (x"02",x"bf",x"6e",x"7e"),
  2393 => (x"4b",x"87",x"c5",x"c0"),
  2394 => (x"0f",x"73",x"49",x"fd"),
  2395 => (x"c1",x"48",x"a6",x"c8"),
  2396 => (x"49",x"fa",x"c3",x"78"),
  2397 => (x"70",x"87",x"e4",x"e0"),
  2398 => (x"02",x"99",x"c2",x"49"),
  2399 => (x"c2",x"87",x"ed",x"c0"),
  2400 => (x"48",x"bf",x"d0",x"f5"),
  2401 => (x"03",x"a8",x"b7",x"c7"),
  2402 => (x"c2",x"87",x"c9",x"c0"),
  2403 => (x"c7",x"48",x"d0",x"f5"),
  2404 => (x"87",x"d3",x"c0",x"78"),
  2405 => (x"c1",x"48",x"66",x"c4"),
  2406 => (x"7e",x"70",x"80",x"e0"),
  2407 => (x"c0",x"02",x"bf",x"6e"),
  2408 => (x"fc",x"4b",x"87",x"c5"),
  2409 => (x"c8",x"0f",x"73",x"49"),
  2410 => (x"78",x"c1",x"48",x"a6"),
  2411 => (x"f5",x"c2",x"7e",x"c0"),
  2412 => (x"50",x"c0",x"48",x"c8"),
  2413 => (x"c3",x"49",x"ee",x"cb"),
  2414 => (x"a6",x"d4",x"87",x"c6"),
  2415 => (x"c8",x"f5",x"c2",x"58"),
  2416 => (x"c1",x"05",x"bf",x"97"),
  2417 => (x"49",x"74",x"87",x"de"),
  2418 => (x"05",x"99",x"f0",x"c3"),
  2419 => (x"c1",x"87",x"cd",x"c0"),
  2420 => (x"df",x"ff",x"49",x"da"),
  2421 => (x"98",x"70",x"87",x"c5"),
  2422 => (x"87",x"c8",x"c1",x"02"),
  2423 => (x"bf",x"e8",x"7e",x"c1"),
  2424 => (x"ff",x"c3",x"49",x"4b"),
  2425 => (x"2b",x"b7",x"c8",x"99"),
  2426 => (x"d9",x"c2",x"b3",x"71"),
  2427 => (x"ff",x"49",x"bf",x"fc"),
  2428 => (x"d0",x"87",x"e6",x"da"),
  2429 => (x"d3",x"c2",x"49",x"66"),
  2430 => (x"02",x"98",x"70",x"87"),
  2431 => (x"c2",x"87",x"c6",x"c0"),
  2432 => (x"c1",x"48",x"c8",x"f5"),
  2433 => (x"c8",x"f5",x"c2",x"50"),
  2434 => (x"c0",x"05",x"bf",x"97"),
  2435 => (x"49",x"73",x"87",x"d6"),
  2436 => (x"05",x"99",x"f0",x"c3"),
  2437 => (x"c1",x"87",x"c5",x"ff"),
  2438 => (x"dd",x"ff",x"49",x"da"),
  2439 => (x"98",x"70",x"87",x"fd"),
  2440 => (x"87",x"f8",x"fe",x"05"),
  2441 => (x"e0",x"c0",x"02",x"6e"),
  2442 => (x"48",x"a6",x"cc",x"87"),
  2443 => (x"bf",x"d0",x"f5",x"c2"),
  2444 => (x"49",x"66",x"cc",x"78"),
  2445 => (x"66",x"c4",x"91",x"cc"),
  2446 => (x"70",x"80",x"71",x"48"),
  2447 => (x"02",x"bf",x"6e",x"7e"),
  2448 => (x"4b",x"87",x"c6",x"c0"),
  2449 => (x"73",x"49",x"66",x"cc"),
  2450 => (x"02",x"66",x"c8",x"0f"),
  2451 => (x"c2",x"87",x"c8",x"c0"),
  2452 => (x"49",x"bf",x"d0",x"f5"),
  2453 => (x"ec",x"87",x"e9",x"f1"),
  2454 => (x"26",x"4d",x"26",x"8e"),
  2455 => (x"26",x"4b",x"26",x"4c"),
  2456 => (x"00",x"00",x"00",x"4f"),
  2457 => (x"00",x"00",x"00",x"00"),
  2458 => (x"14",x"11",x"12",x"58"),
  2459 => (x"23",x"1c",x"1b",x"1d"),
  2460 => (x"94",x"91",x"59",x"5a"),
  2461 => (x"f4",x"eb",x"f2",x"f5"),
  2462 => (x"00",x"00",x"00",x"00"),
  2463 => (x"00",x"00",x"00",x"00"),
  2464 => (x"ff",x"4a",x"71",x"1e"),
  2465 => (x"72",x"49",x"bf",x"c8"),
  2466 => (x"4f",x"26",x"48",x"a1"),
  2467 => (x"bf",x"c8",x"ff",x"1e"),
  2468 => (x"c0",x"c0",x"fe",x"89"),
  2469 => (x"a9",x"c0",x"c0",x"c0"),
  2470 => (x"c0",x"87",x"c4",x"01"),
  2471 => (x"c1",x"87",x"c2",x"4a"),
  2472 => (x"26",x"48",x"72",x"4a"),
  2473 => (x"5b",x"5e",x"0e",x"4f"),
  2474 => (x"71",x"0e",x"5d",x"5c"),
  2475 => (x"4c",x"d4",x"ff",x"4b"),
  2476 => (x"c0",x"48",x"66",x"d0"),
  2477 => (x"ff",x"49",x"d6",x"78"),
  2478 => (x"c3",x"87",x"dd",x"dd"),
  2479 => (x"49",x"6c",x"7c",x"ff"),
  2480 => (x"71",x"99",x"ff",x"c3"),
  2481 => (x"f0",x"c3",x"49",x"4d"),
  2482 => (x"a9",x"e0",x"c1",x"99"),
  2483 => (x"c3",x"87",x"cb",x"05"),
  2484 => (x"48",x"6c",x"7c",x"ff"),
  2485 => (x"66",x"d0",x"98",x"c3"),
  2486 => (x"ff",x"c3",x"78",x"08"),
  2487 => (x"49",x"4a",x"6c",x"7c"),
  2488 => (x"ff",x"c3",x"31",x"c8"),
  2489 => (x"71",x"4a",x"6c",x"7c"),
  2490 => (x"c8",x"49",x"72",x"b2"),
  2491 => (x"7c",x"ff",x"c3",x"31"),
  2492 => (x"b2",x"71",x"4a",x"6c"),
  2493 => (x"31",x"c8",x"49",x"72"),
  2494 => (x"6c",x"7c",x"ff",x"c3"),
  2495 => (x"ff",x"b2",x"71",x"4a"),
  2496 => (x"e0",x"c0",x"48",x"d0"),
  2497 => (x"02",x"9b",x"73",x"78"),
  2498 => (x"7b",x"72",x"87",x"c2"),
  2499 => (x"4d",x"26",x"48",x"75"),
  2500 => (x"4b",x"26",x"4c",x"26"),
  2501 => (x"26",x"1e",x"4f",x"26"),
  2502 => (x"5b",x"5e",x"0e",x"4f"),
  2503 => (x"86",x"f8",x"0e",x"5c"),
  2504 => (x"a6",x"c8",x"1e",x"76"),
  2505 => (x"87",x"fd",x"fd",x"49"),
  2506 => (x"4b",x"70",x"86",x"c4"),
  2507 => (x"a8",x"c2",x"48",x"6e"),
  2508 => (x"87",x"f0",x"c2",x"03"),
  2509 => (x"f0",x"c3",x"4a",x"73"),
  2510 => (x"aa",x"d0",x"c1",x"9a"),
  2511 => (x"c1",x"87",x"c7",x"02"),
  2512 => (x"c2",x"05",x"aa",x"e0"),
  2513 => (x"49",x"73",x"87",x"de"),
  2514 => (x"c3",x"02",x"99",x"c8"),
  2515 => (x"87",x"c6",x"ff",x"87"),
  2516 => (x"9c",x"c3",x"4c",x"73"),
  2517 => (x"c1",x"05",x"ac",x"c2"),
  2518 => (x"66",x"c4",x"87",x"c2"),
  2519 => (x"71",x"31",x"c9",x"49"),
  2520 => (x"4a",x"66",x"c4",x"1e"),
  2521 => (x"f5",x"c2",x"92",x"d4"),
  2522 => (x"81",x"72",x"49",x"d4"),
  2523 => (x"87",x"e4",x"cd",x"fe"),
  2524 => (x"da",x"ff",x"49",x"d8"),
  2525 => (x"c0",x"c8",x"87",x"e2"),
  2526 => (x"ec",x"e3",x"c2",x"1e"),
  2527 => (x"d6",x"e7",x"fd",x"49"),
  2528 => (x"48",x"d0",x"ff",x"87"),
  2529 => (x"c2",x"78",x"e0",x"c0"),
  2530 => (x"cc",x"1e",x"ec",x"e3"),
  2531 => (x"92",x"d4",x"4a",x"66"),
  2532 => (x"49",x"d4",x"f5",x"c2"),
  2533 => (x"cb",x"fe",x"81",x"72"),
  2534 => (x"86",x"cc",x"87",x"eb"),
  2535 => (x"c1",x"05",x"ac",x"c1"),
  2536 => (x"66",x"c4",x"87",x"c2"),
  2537 => (x"71",x"31",x"c9",x"49"),
  2538 => (x"4a",x"66",x"c4",x"1e"),
  2539 => (x"f5",x"c2",x"92",x"d4"),
  2540 => (x"81",x"72",x"49",x"d4"),
  2541 => (x"87",x"dc",x"cc",x"fe"),
  2542 => (x"1e",x"ec",x"e3",x"c2"),
  2543 => (x"d4",x"4a",x"66",x"c8"),
  2544 => (x"d4",x"f5",x"c2",x"92"),
  2545 => (x"fe",x"81",x"72",x"49"),
  2546 => (x"d7",x"87",x"eb",x"c9"),
  2547 => (x"c7",x"d9",x"ff",x"49"),
  2548 => (x"1e",x"c0",x"c8",x"87"),
  2549 => (x"49",x"ec",x"e3",x"c2"),
  2550 => (x"87",x"d8",x"e5",x"fd"),
  2551 => (x"d0",x"ff",x"86",x"cc"),
  2552 => (x"78",x"e0",x"c0",x"48"),
  2553 => (x"4c",x"26",x"8e",x"f8"),
  2554 => (x"4f",x"26",x"4b",x"26"),
  2555 => (x"5c",x"5b",x"5e",x"0e"),
  2556 => (x"86",x"fc",x"0e",x"5d"),
  2557 => (x"d4",x"ff",x"4d",x"71"),
  2558 => (x"7e",x"66",x"d4",x"4c"),
  2559 => (x"a8",x"b7",x"c3",x"48"),
  2560 => (x"87",x"e2",x"c1",x"01"),
  2561 => (x"66",x"c4",x"1e",x"75"),
  2562 => (x"c2",x"93",x"d4",x"4b"),
  2563 => (x"73",x"83",x"d4",x"f5"),
  2564 => (x"e0",x"c3",x"fe",x"49"),
  2565 => (x"49",x"a3",x"c8",x"87"),
  2566 => (x"d0",x"ff",x"49",x"69"),
  2567 => (x"78",x"e1",x"c8",x"48"),
  2568 => (x"48",x"71",x"7c",x"dd"),
  2569 => (x"70",x"98",x"ff",x"c3"),
  2570 => (x"c8",x"4a",x"71",x"7c"),
  2571 => (x"48",x"72",x"2a",x"b7"),
  2572 => (x"70",x"98",x"ff",x"c3"),
  2573 => (x"d0",x"4a",x"71",x"7c"),
  2574 => (x"48",x"72",x"2a",x"b7"),
  2575 => (x"70",x"98",x"ff",x"c3"),
  2576 => (x"d8",x"48",x"71",x"7c"),
  2577 => (x"7c",x"70",x"28",x"b7"),
  2578 => (x"7c",x"7c",x"7c",x"c0"),
  2579 => (x"7c",x"7c",x"7c",x"7c"),
  2580 => (x"7c",x"7c",x"7c",x"7c"),
  2581 => (x"48",x"d0",x"ff",x"7c"),
  2582 => (x"c4",x"78",x"e0",x"c0"),
  2583 => (x"49",x"dc",x"1e",x"66"),
  2584 => (x"87",x"d9",x"d7",x"ff"),
  2585 => (x"8e",x"fc",x"86",x"c8"),
  2586 => (x"4c",x"26",x"4d",x"26"),
  2587 => (x"4f",x"26",x"4b",x"26"),
  2588 => (x"c0",x"1e",x"73",x"1e"),
  2589 => (x"f0",x"e2",x"c2",x"4b"),
  2590 => (x"c2",x"50",x"c0",x"48"),
  2591 => (x"49",x"bf",x"ec",x"e2"),
  2592 => (x"87",x"c2",x"dc",x"fe"),
  2593 => (x"c4",x"05",x"98",x"70"),
  2594 => (x"d4",x"e2",x"c2",x"87"),
  2595 => (x"26",x"48",x"73",x"4b"),
  2596 => (x"00",x"4f",x"26",x"4b"),
  2597 => (x"77",x"6f",x"68",x"53"),
  2598 => (x"64",x"69",x"68",x"2f"),
  2599 => (x"53",x"4f",x"20",x"65"),
  2600 => (x"20",x"3d",x"20",x"44"),
  2601 => (x"20",x"79",x"65",x"6b"),
  2602 => (x"00",x"32",x"31",x"46"),
  2603 => (x"00",x"00",x"28",x"b4"),
  2604 => (x"00",x"00",x"00",x"00"),
  2605 => (x"4f",x"54",x"55",x"41"),
  2606 => (x"54",x"4f",x"4f",x"42"),
  2607 => (x"00",x"53",x"45",x"4e"),
  2608 => (x"00",x"00",x"1b",x"af"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

